module adder_i52_o27 (a,b,r);
input [25:0] a,b;
output [26:0] r;

assign r = a+b;

endmodule

