module adder_i24_o13 (a,b,r);
input [11:0] a,b;
output [12:0] r;

assign r = a+b;

endmodule

