module adder_i56_o29 (a,b,r);
input [27:0] a,b;
output [28:0] r;

assign r = a+b;

endmodule

