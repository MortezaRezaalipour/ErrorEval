module top(pi0, pi1, pi2, pi3, pi4, pi5, po0, po1, po2, po3);
  input pi0, pi1, pi2, pi3, pi4, pi5;
  output po0, po1, po2, po3;
  wire n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27;
  assign n7 = pi0 & pi2;
  assign n8 = pi4 & n7;
  assign n9 = ~pi4 & ~n7;
  assign n10 = ~n8 & ~n9;
  assign n11 = pi0 & pi3;
  assign n12 = pi1 & pi2;
  assign n13 = pi5 & n12;
  assign n14 = ~pi5 & ~n12;
  assign n15 = ~n13 & ~n14;
  assign n16 = n11 & n15;
  assign n17 = ~n11 & ~n15;
  assign n18 = ~n16 & ~n17;
  assign n19 = n8 & n18;
  assign n20 = ~n8 & ~n18;
  assign n21 = ~n19 & ~n20;
  assign n22 = pi1 & pi3;
  assign n23 = ~n13 & ~n16;
  assign n24 = n22 & ~n23;
  assign n25 = ~n22 & n23;
  assign n26 = ~n24 & ~n25;
  assign n27 = ~n19 & ~n26;
  assign po0 = n10;
  assign po1 = n21;
  assign po2 = ~n27;
  assign po3 = n24;
endmodule
