module multiplier (a, b, r);
input [1:0] a, b;
output [2:0] r;


assign r = a * b;

endmodule 
