// Benchmark "circuit" written by ABC on Tue Apr 12 03:26:52 2022

module circuit ( 
    g0, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11,
    g378, g377, g376, g375, g374, g373, g372, g371, g370, g369, g368, g367  );
  input  g0, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11;
  output g378, g377, g376, g375, g374, g373, g372, g371, g370, g369, g368,
    g367;
  wire g12, g13, g14, g15, g16, g17, g18, g19, g20, g21, g22, g23, g24, g25,
    g26, g27, g28, g29, g30, g31, g32, g33, g34, g35, g36, g37, g38, g39,
    g40, g41, g42, g43, g44, g45, g46, g47, g48, g49, g50, g51, g52, g53,
    g54, g55, g56, g57, g58, g59, g60, g61, g62, g63, g64, g65, g66, g67,
    g68, g69, g70, g71, g72, g73, g74, g75, g76, g77, g78, g79, g80, g81,
    g82, g83, g84, g85, g86, g87, g88, g89, g90, g91, g92, g93, g94, g95,
    g96, g97, g98, g99, g100, g101, g102, g103, g104, g105, g106, g107,
    g108, g109, g110, g111, g112, g113, g114, g115, g116, g117, g118, g119,
    g120, g121, g122, g123, g124, g125, g126, g127, g128, g129, g130, g131,
    g132, g133, g134, g135, g136, g137, g138, g139, g140, g141, g142, g143,
    g144, g145, g146, g147, g148, g149, g150, g151, g152, g153, g154, g155,
    g156, g157, g158, g159, g160, g161, g162, g163, g164, g165, g166, g167,
    g168, g169, g170, g171, g172, g173, g174, g175, g176, g177, g178, g179,
    g180, g181, g182, g183, g184, g185, g186, g187, g188, g189, g190, g191,
    g192, g193, g194, g195, g196, g197, g198, g199, g200, g201, g202, g203,
    g204, g205, g206, g207, g208, g209, g210, g211, g212, g213, g214, g215,
    g216, g217, g218, g219, g220, g221, g222, g223, g224, g225, g226, g227,
    g228, g229, g230, g231, g232, g233, g234, g235, g236, g237, g238, g239,
    g240, g241, g242, g243, g244, g245, g246, g247, g248, g249, g250, g251,
    g252, g253, g254, g255, g256, g257, g258, g259, g260, g261, g262, g263,
    g264, g265, g266, g267, g268, g269, g270, g271, g272, g273, g274, g275,
    g276, g277, g278, g279, g280, g281, g282, g283, g284, g285, g286, g287,
    g288, g289, g290, g291, g292, g293, g294, g295, g296, g297, g298, g299,
    g300, g301, g302, g303, g304, g305, g306, g307, g308, g309, g310, g311,
    g312, g313, g314, g315, g316, g317, g318, g319, g320, g321, g322, g323,
    g324, g325, g326, g327, g328, g329, g330, g331, g332, g333, g334, g335,
    g336, g337, g338, g339, g340, g341, g342, g343, g344, g345, g346, g347,
    g348, g349, g350, g351, g352, g353, g354, g355, g356, g357, g358, g359,
    g360, g361, g362, g363, g364, g365, g366;
  assign g12 = 1'b0;
  assign g13 = 1'b0;
  assign g14 = 1'b0;
  assign g15 = 1'b0;
  assign g16 = 1'b0;
  assign g17 = 1'b0;
  assign g18 = 1'b0;
  assign g19 = 1'b0;
  assign g20 = 1'b0;
  assign g21 = 1'b0;
  assign g22 = 1'b0;
  assign g23 = 1'b0;
  assign g24 = 1'b0;
  assign g25 = 1'b0;
  assign g26 = 1'b0;
  assign g27 = 1'b0;
  assign g28 = 1'b0;
  assign g29 = 1'b0;
  assign g30 = 1'b0;
  assign g31 = 1'b0;
  assign g32 = 1'b0;
  assign g33 = 1'b0;
  assign g34 = 1'b0;
  assign g35 = g4 & g8;
  assign g36 = 1'b0;
  assign g37 = 1'b0;
  assign g38 = 1'b0;
  assign g39 = 1'b0;
  assign g40 = 1'b0;
  assign g41 = 1'b0;
  assign g42 = 1'b0;
  assign g43 = 1'b0;
  assign g44 = 1'b0;
  assign g45 = 1'b0;
  assign g46 = 1'b0;
  assign g47 = 1'b0;
  assign g48 = 1'b0;
  assign g49 = 1'b0;
  assign g50 = 1'b0;
  assign g51 = 1'b0;
  assign g52 = 1'b0;
  assign g53 = 1'b0;
  assign g54 = 1'b0;
  assign g55 = 1'b0;
  assign g56 = 1'b0;
  assign g57 = 1'b0;
  assign g58 = 1'b0;
  assign g59 = 1'b0;
  assign g60 = 1'b0;
  assign g61 = 1'b0;
  assign g62 = 1'b0;
  assign g63 = 1'b0;
  assign g64 = 1'b0;
  assign g65 = 1'b0;
  assign g66 = 1'b0;
  assign g67 = 1'b0;
  assign g68 = 1'b0;
  assign g69 = 1'b0;
  assign g70 = 1'b0;
  assign g71 = 1'b0;
  assign g72 = 1'b0;
  assign g73 = 1'b0;
  assign g74 = 1'b0;
  assign g75 = 1'b0;
  assign g76 = 1'b0;
  assign g77 = 1'b0;
  assign g78 = 1'b0;
  assign g79 = 1'b0;
  assign g80 = 1'b0;
  assign g81 = 1'b0;
  assign g82 = 1'b0;
  assign g83 = 1'b0;
  assign g84 = 1'b0;
  assign g85 = 1'b0;
  assign g86 = 1'b0;
  assign g87 = 1'b0;
  assign g88 = 1'b0;
  assign g89 = 1'b0;
  assign g90 = 1'b0;
  assign g91 = 1'b0;
  assign g92 = 1'b0;
  assign g93 = 1'b0;
  assign g94 = 1'b0;
  assign g95 = 1'b0;
  assign g96 = 1'b0;
  assign g97 = 1'b0;
  assign g98 = 1'b0;
  assign g99 = 1'b0;
  assign g100 = 1'b0;
  assign g101 = 1'b0;
  assign g102 = 1'b0;
  assign g103 = 1'b0;
  assign g104 = 1'b0;
  assign g105 = 1'b0;
  assign g106 = 1'b0;
  assign g107 = 1'b0;
  assign g108 = 1'b0;
  assign g109 = 1'b0;
  assign g110 = 1'b0;
  assign g111 = 1'b0;
  assign g112 = 1'b0;
  assign g113 = 1'b0;
  assign g114 = 1'b0;
  assign g115 = 1'b0;
  assign g116 = 1'b0;
  assign g117 = 1'b0;
  assign g118 = 1'b0;
  assign g119 = 1'b0;
  assign g120 = 1'b0;
  assign g121 = 1'b0;
  assign g122 = 1'b0;
  assign g123 = 1'b0;
  assign g124 = 1'b0;
  assign g125 = 1'b0;
  assign g126 = 1'b0;
  assign g127 = 1'b0;
  assign g128 = 1'b0;
  assign g129 = 1'b0;
  assign g130 = 1'b0;
  assign g131 = 1'b0;
  assign g132 = 1'b0;
  assign g133 = 1'b0;
  assign g134 = 1'b0;
  assign g135 = 1'b0;
  assign g136 = 1'b0;
  assign g137 = 1'b0;
  assign g138 = 1'b0;
  assign g139 = 1'b0;
  assign g140 = 1'b0;
  assign g141 = 1'b0;
  assign g142 = 1'b0;
  assign g143 = 1'b0;
  assign g144 = 1'b0;
  assign g145 = 1'b0;
  assign g146 = 1'b0;
  assign g147 = 1'b0;
  assign g148 = 1'b0;
  assign g149 = 1'b0;
  assign g150 = 1'b0;
  assign g151 = 1'b0;
  assign g152 = 1'b0;
  assign g153 = 1'b0;
  assign g154 = 1'b0;
  assign g155 = 1'b0;
  assign g156 = 1'b0;
  assign g157 = 1'b0;
  assign g158 = 1'b0;
  assign g159 = 1'b0;
  assign g160 = 1'b0;
  assign g161 = 1'b0;
  assign g162 = 1'b0;
  assign g163 = 1'b0;
  assign g164 = 1'b0;
  assign g165 = 1'b0;
  assign g166 = 1'b0;
  assign g167 = 1'b0;
  assign g168 = 1'b0;
  assign g169 = 1'b0;
  assign g170 = 1'b0;
  assign g171 = 1'b0;
  assign g172 = 1'b0;
  assign g173 = 1'b0;
  assign g174 = 1'b0;
  assign g175 = 1'b0;
  assign g176 = 1'b0;
  assign g177 = 1'b0;
  assign g178 = 1'b0;
  assign g179 = 1'b0;
  assign g180 = 1'b0;
  assign g181 = 1'b0;
  assign g182 = 1'b0;
  assign g183 = 1'b0;
  assign g184 = 1'b0;
  assign g185 = 1'b0;
  assign g186 = 1'b0;
  assign g187 = 1'b0;
  assign g188 = 1'b0;
  assign g189 = 1'b0;
  assign g190 = 1'b0;
  assign g191 = 1'b0;
  assign g192 = 1'b0;
  assign g193 = 1'b0;
  assign g194 = 1'b0;
  assign g195 = 1'b0;
  assign g196 = 1'b0;
  assign g197 = 1'b0;
  assign g198 = 1'b0;
  assign g199 = 1'b0;
  assign g200 = 1'b0;
  assign g201 = 1'b0;
  assign g202 = 1'b0;
  assign g203 = 1'b0;
  assign g204 = 1'b0;
  assign g205 = 1'b0;
  assign g206 = 1'b0;
  assign g207 = 1'b0;
  assign g208 = 1'b0;
  assign g209 = 1'b0;
  assign g210 = 1'b0;
  assign g211 = 1'b0;
  assign g212 = 1'b0;
  assign g213 = 1'b0;
  assign g214 = 1'b0;
  assign g215 = 1'b0;
  assign g216 = 1'b0;
  assign g217 = 1'b0;
  assign g218 = 1'b0;
  assign g219 = 1'b0;
  assign g220 = 1'b0;
  assign g221 = 1'b0;
  assign g222 = 1'b0;
  assign g223 = 1'b0;
  assign g224 = 1'b0;
  assign g225 = 1'b0;
  assign g226 = 1'b0;
  assign g227 = 1'b0;
  assign g228 = 1'b0;
  assign g229 = 1'b0;
  assign g230 = 1'b0;
  assign g231 = 1'b0;
  assign g232 = 1'b0;
  assign g233 = 1'b0;
  assign g234 = 1'b0;
  assign g235 = 1'b0;
  assign g236 = 1'b0;
  assign g237 = 1'b0;
  assign g238 = 1'b0;
  assign g239 = 1'b0;
  assign g240 = 1'b0;
  assign g241 = 1'b0;
  assign g242 = 1'b0;
  assign g243 = 1'b0;
  assign g244 = 1'b0;
  assign g245 = 1'b0;
  assign g246 = 1'b0;
  assign g247 = 1'b0;
  assign g248 = 1'b0;
  assign g249 = 1'b0;
  assign g250 = 1'b0;
  assign g251 = 1'b0;
  assign g252 = 1'b0;
  assign g253 = 1'b0;
  assign g254 = 1'b0;
  assign g255 = 1'b0;
  assign g256 = 1'b0;
  assign g257 = 1'b0;
  assign g258 = 1'b0;
  assign g259 = 1'b0;
  assign g260 = 1'b0;
  assign g261 = 1'b0;
  assign g262 = 1'b0;
  assign g263 = 1'b0;
  assign g264 = 1'b0;
  assign g265 = 1'b0;
  assign g266 = 1'b0;
  assign g267 = 1'b0;
  assign g268 = 1'b0;
  assign g269 = 1'b0;
  assign g270 = 1'b0;
  assign g271 = 1'b0;
  assign g272 = 1'b0;
  assign g273 = 1'b0;
  assign g274 = 1'b0;
  assign g275 = 1'b0;
  assign g276 = 1'b0;
  assign g277 = 1'b0;
  assign g278 = 1'b0;
  assign g279 = 1'b0;
  assign g280 = 1'b0;
  assign g281 = 1'b0;
  assign g282 = 1'b0;
  assign g283 = 1'b0;
  assign g284 = 1'b0;
  assign g285 = 1'b0;
  assign g286 = 1'b0;
  assign g287 = 1'b0;
  assign g288 = 1'b0;
  assign g289 = 1'b0;
  assign g290 = 1'b0;
  assign g291 = 1'b0;
  assign g292 = 1'b0;
  assign g293 = 1'b0;
  assign g294 = 1'b0;
  assign g295 = 1'b0;
  assign g296 = 1'b0;
  assign g297 = 1'b0;
  assign g298 = 1'b0;
  assign g299 = 1'b0;
  assign g300 = 1'b0;
  assign g301 = 1'b0;
  assign g302 = 1'b0;
  assign g303 = 1'b0;
  assign g304 = 1'b0;
  assign g305 = 1'b0;
  assign g306 = 1'b0;
  assign g307 = 1'b0;
  assign g308 = 1'b0;
  assign g309 = 1'b0;
  assign g310 = 1'b0;
  assign g311 = 1'b0;
  assign g312 = 1'b0;
  assign g313 = 1'b0;
  assign g314 = 1'b0;
  assign g315 = 1'b0;
  assign g316 = 1'b0;
  assign g317 = 1'b0;
  assign g318 = 1'b0;
  assign g319 = 1'b0;
  assign g320 = 1'b0;
  assign g321 = 1'b0;
  assign g322 = 1'b0;
  assign g323 = 1'b0;
  assign g324 = 1'b0;
  assign g325 = 1'b0;
  assign g326 = 1'b0;
  assign g327 = 1'b0;
  assign g328 = 1'b0;
  assign g329 = 1'b0;
  assign g330 = 1'b0;
  assign g331 = 1'b0;
  assign g332 = 1'b0;
  assign g333 = 1'b0;
  assign g334 = 1'b0;
  assign g335 = 1'b0;
  assign g336 = 1'b0;
  assign g337 = 1'b0;
  assign g338 = 1'b0;
  assign g339 = 1'b0;
  assign g340 = 1'b0;
  assign g341 = 1'b0;
  assign g342 = 1'b0;
  assign g343 = 1'b0;
  assign g344 = 1'b0;
  assign g345 = 1'b0;
  assign g346 = 1'b0;
  assign g347 = 1'b0;
  assign g348 = 1'b0;
  assign g349 = 1'b0;
  assign g350 = 1'b0;
  assign g351 = 1'b0;
  assign g352 = 1'b0;
  assign g353 = 1'b0;
  assign g354 = 1'b0;
  assign g355 = 1'b0;
  assign g356 = 1'b0;
  assign g357 = 1'b0;
  assign g358 = 1'b0;
  assign g359 = 1'b0;
  assign g360 = 1'b0;
  assign g361 = 1'b0;
  assign g362 = 1'b0;
  assign g363 = 1'b0;
  assign g364 = 1'b0;
  assign g365 = 1'b0;
  assign g366 = 1'b0;
  assign g367 = g366;
  assign g368 = g187;
  assign g369 = g203;
  assign g370 = g231;
  assign g371 = g266;
  assign g372 = g295;
  assign g373 = g317;
  assign g374 = g339;
  assign g375 = g352;
  assign g376 = g358;
  assign g377 = g365;
  assign g378 = g363;
endmodule


