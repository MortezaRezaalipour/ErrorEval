module madd_8_app2(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15;
  wire n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538;
  assign n25 = pi02 & pi09;
  assign n26 = pi03 & pi10;
  assign n27 = n25 & n26;
  assign n28 = pi05 & pi08;
  assign n29 = n27 & n28;
  assign n30 = ~n27 & ~n28;
  assign n31 = ~n29 & ~n30;
  assign n32 = pi04 & pi09;
  assign n33 = n26 & n32;
  assign n34 = ~n26 & ~n32;
  assign n35 = ~n33 & ~n34;
  assign n36 = n31 & n35;
  assign n37 = ~n29 & ~n36;
  assign n38 = pi01 & pi12;
  assign n39 = pi00 & pi13;
  assign n40 = n38 & n39;
  assign n41 = pi02 & pi11;
  assign n42 = ~n38 & ~n39;
  assign n43 = ~n40 & ~n42;
  assign n44 = n41 & n43;
  assign n45 = ~n40 & ~n44;
  assign n46 = pi05 & pi10;
  assign n47 = n32 & n46;
  assign n48 = pi04 & pi10;
  assign n49 = pi05 & pi09;
  assign n50 = ~n48 & ~n49;
  assign n51 = ~n47 & ~n50;
  assign n52 = ~n45 & n51;
  assign n53 = n45 & ~n51;
  assign n54 = ~n52 & ~n53;
  assign n55 = ~n37 & n54;
  assign n56 = n37 & ~n54;
  assign n57 = ~n55 & ~n56;
  assign n58 = pi01 & pi14;
  assign n59 = n39 & n58;
  assign n60 = pi01 & pi13;
  assign n61 = pi00 & pi14;
  assign n62 = ~n60 & ~n61;
  assign n63 = ~n59 & ~n62;
  assign n64 = pi06 & pi08;
  assign n65 = ~n63 & ~n64;
  assign n66 = n63 & n64;
  assign n67 = ~n65 & ~n66;
  assign n68 = pi03 & pi12;
  assign n69 = n41 & n68;
  assign n70 = pi02 & pi12;
  assign n71 = pi03 & pi11;
  assign n72 = ~n70 & ~n71;
  assign n73 = ~n69 & ~n72;
  assign n74 = n33 & n73;
  assign n75 = ~n33 & ~n73;
  assign n76 = ~n74 & ~n75;
  assign n77 = ~n67 & ~n76;
  assign n78 = n67 & n76;
  assign n79 = ~n77 & ~n78;
  assign n80 = ~n41 & ~n43;
  assign n81 = ~n44 & ~n80;
  assign n82 = pi00 & pi11;
  assign n83 = n38 & n82;
  assign n84 = pi00 & pi12;
  assign n85 = pi01 & pi11;
  assign n86 = ~n84 & ~n85;
  assign n87 = ~n83 & ~n86;
  assign n88 = pi04 & pi08;
  assign n89 = n87 & n88;
  assign n90 = ~n83 & ~n89;
  assign n91 = n81 & ~n90;
  assign n92 = ~n81 & n90;
  assign n93 = ~n91 & ~n92;
  assign n94 = pi00 & pi09;
  assign n95 = n41 & n94;
  assign n96 = pi02 & pi10;
  assign n97 = pi03 & pi09;
  assign n98 = ~n96 & ~n97;
  assign n99 = ~n27 & ~n98;
  assign n100 = n95 & n99;
  assign n101 = ~n95 & ~n99;
  assign n102 = ~n100 & ~n101;
  assign n103 = pi01 & pi10;
  assign n104 = n94 & n103;
  assign n105 = pi03 & pi08;
  assign n106 = n103 & n105;
  assign n107 = ~n104 & ~n106;
  assign n108 = n102 & ~n107;
  assign n109 = ~n100 & ~n108;
  assign n110 = n93 & ~n109;
  assign n111 = ~n91 & ~n110;
  assign n112 = n79 & ~n111;
  assign n113 = ~n79 & n111;
  assign n114 = ~n112 & ~n113;
  assign n115 = n57 & n114;
  assign n116 = ~n57 & ~n114;
  assign n117 = ~n115 & ~n116;
  assign n118 = ~n93 & n109;
  assign n119 = ~n110 & ~n118;
  assign n120 = ~n31 & ~n35;
  assign n121 = ~n36 & ~n120;
  assign n122 = n119 & n121;
  assign n123 = ~n119 & ~n121;
  assign n124 = ~n122 & ~n123;
  assign n125 = ~n87 & ~n88;
  assign n126 = ~n89 & ~n125;
  assign n127 = ~n102 & n107;
  assign n128 = ~n108 & ~n127;
  assign n129 = n126 & n128;
  assign n130 = ~n126 & ~n128;
  assign n131 = ~n129 & ~n130;
  assign n132 = ~n25 & ~n82;
  assign n133 = ~n95 & ~n132;
  assign n134 = ~n94 & n103;
  assign n135 = n105 & ~n134;
  assign n136 = ~n105 & n134;
  assign n137 = ~n135 & ~n136;
  assign n138 = n133 & ~n137;
  assign n139 = ~n105 & ~n134;
  assign n140 = n105 & n134;
  assign n141 = ~n139 & ~n140;
  assign n142 = ~n133 & ~n141;
  assign n143 = ~n138 & ~n142;
  assign n144 = pi01 & pi09;
  assign n145 = pi00 & pi10;
  assign n146 = ~n144 & ~n145;
  assign n147 = ~n104 & ~n146;
  assign n148 = pi02 & pi08;
  assign n149 = n147 & n148;
  assign n150 = pi01 & pi08;
  assign n151 = n94 & n150;
  assign n152 = ~n147 & ~n148;
  assign n153 = ~n149 & ~n152;
  assign n154 = n151 & n153;
  assign n155 = ~n149 & ~n154;
  assign n156 = n143 & ~n155;
  assign n157 = ~n138 & ~n156;
  assign n158 = n131 & ~n157;
  assign n159 = ~n129 & ~n158;
  assign n160 = n124 & ~n159;
  assign n161 = ~n122 & ~n160;
  assign n162 = ~n117 & n161;
  assign n163 = n117 & ~n161;
  assign n164 = ~n162 & ~n163;
  assign n165 = ~n151 & ~n153;
  assign n166 = ~n154 & ~n165;
  assign n167 = pi00 & pi08;
  assign n168 = pi16 & n167;
  assign n169 = ~pi17 & ~n168;
  assign n170 = pi17 & n168;
  assign n171 = ~n94 & ~n150;
  assign n172 = ~n151 & ~n171;
  assign n173 = ~n170 & ~n172;
  assign n174 = ~n169 & ~n173;
  assign n175 = ~n166 & ~n174;
  assign n176 = ~n169 & n172;
  assign n177 = ~n170 & ~n176;
  assign n178 = n166 & ~n177;
  assign n179 = ~pi18 & ~n178;
  assign n180 = ~n175 & ~n179;
  assign n181 = ~n143 & n155;
  assign n182 = ~n156 & ~n181;
  assign n183 = ~n180 & ~n182;
  assign n184 = pi18 & ~n175;
  assign n185 = ~n178 & ~n184;
  assign n186 = n182 & ~n185;
  assign n187 = ~pi19 & ~n186;
  assign n188 = ~n183 & ~n187;
  assign n189 = ~n131 & n157;
  assign n190 = ~n158 & ~n189;
  assign n191 = ~n188 & ~n190;
  assign n192 = pi19 & ~n183;
  assign n193 = ~n186 & ~n192;
  assign n194 = n190 & ~n193;
  assign n195 = ~pi20 & ~n194;
  assign n196 = ~n191 & ~n195;
  assign n197 = ~n124 & n159;
  assign n198 = ~n160 & ~n197;
  assign n199 = n196 & n198;
  assign n200 = ~n196 & ~n198;
  assign n201 = pi21 & ~n200;
  assign n202 = ~n199 & ~n201;
  assign n203 = n164 & ~n202;
  assign n204 = ~n164 & n202;
  assign n205 = pi22 & ~n204;
  assign n206 = ~n203 & ~n205;
  assign n207 = ~n52 & ~n55;
  assign n208 = ~n59 & ~n66;
  assign n209 = pi06 & pi09;
  assign n210 = ~n32 & n46;
  assign n211 = n209 & ~n210;
  assign n212 = ~n209 & n210;
  assign n213 = ~n211 & ~n212;
  assign n214 = ~n208 & ~n213;
  assign n215 = ~n209 & ~n210;
  assign n216 = n209 & n210;
  assign n217 = ~n215 & ~n216;
  assign n218 = n208 & ~n217;
  assign n219 = ~n214 & ~n218;
  assign n220 = ~n207 & n219;
  assign n221 = n207 & ~n219;
  assign n222 = ~n220 & ~n221;
  assign n223 = ~n78 & ~n112;
  assign n224 = ~n222 & n223;
  assign n225 = n222 & ~n223;
  assign n226 = ~n224 & ~n225;
  assign n227 = pi00 & pi15;
  assign n228 = n58 & n227;
  assign n229 = ~n58 & ~n227;
  assign n230 = ~n228 & ~n229;
  assign n231 = pi04 & pi11;
  assign n232 = ~n230 & ~n231;
  assign n233 = n230 & n231;
  assign n234 = ~n232 & ~n233;
  assign n235 = ~n69 & ~n74;
  assign n236 = pi02 & pi13;
  assign n237 = pi07 & pi12;
  assign n238 = n105 & n237;
  assign n239 = pi07 & pi08;
  assign n240 = ~n68 & ~n239;
  assign n241 = ~n238 & ~n240;
  assign n242 = n236 & n241;
  assign n243 = ~n236 & ~n241;
  assign n244 = ~n242 & ~n243;
  assign n245 = ~n235 & n244;
  assign n246 = n235 & ~n244;
  assign n247 = ~n245 & ~n246;
  assign n248 = n234 & n247;
  assign n249 = ~n234 & ~n247;
  assign n250 = ~n248 & ~n249;
  assign n251 = ~n226 & ~n250;
  assign n252 = n226 & n250;
  assign n253 = ~n251 & ~n252;
  assign n254 = ~n115 & ~n163;
  assign n255 = n253 & ~n254;
  assign n256 = ~n253 & n254;
  assign n257 = ~n255 & ~n256;
  assign n258 = ~n206 & n257;
  assign n259 = ~pi22 & ~n203;
  assign n260 = ~n204 & ~n259;
  assign n261 = ~n257 & ~n260;
  assign n262 = pi23 & ~n261;
  assign n263 = ~n258 & ~n262;
  assign n264 = ~n252 & ~n255;
  assign n265 = ~pi06 & n47;
  assign n266 = ~n214 & ~n265;
  assign n267 = n46 & n209;
  assign n268 = pi03 & pi14;
  assign n269 = n236 & n268;
  assign n270 = pi02 & pi14;
  assign n271 = pi03 & pi13;
  assign n272 = ~n270 & ~n271;
  assign n273 = ~n269 & ~n272;
  assign n274 = ~n267 & ~n273;
  assign n275 = n267 & n273;
  assign n276 = ~n274 & ~n275;
  assign n277 = pi04 & pi12;
  assign n278 = pi05 & pi11;
  assign n279 = n277 & n278;
  assign n280 = ~n277 & ~n278;
  assign n281 = ~n279 & ~n280;
  assign n282 = pi07 & pi09;
  assign n283 = n281 & n282;
  assign n284 = ~n281 & ~n282;
  assign n285 = ~n283 & ~n284;
  assign n286 = ~n276 & ~n285;
  assign n287 = n276 & n285;
  assign n288 = ~n286 & ~n287;
  assign n289 = ~n266 & n288;
  assign n290 = n266 & ~n288;
  assign n291 = ~n289 & ~n290;
  assign n292 = ~n245 & ~n248;
  assign n293 = ~n238 & ~n242;
  assign n294 = ~n228 & ~n233;
  assign n295 = pi06 & pi15;
  assign n296 = n103 & n295;
  assign n297 = pi01 & pi15;
  assign n298 = pi06 & pi10;
  assign n299 = ~n297 & ~n298;
  assign n300 = ~n296 & ~n299;
  assign n301 = ~n294 & n300;
  assign n302 = n294 & ~n300;
  assign n303 = ~n301 & ~n302;
  assign n304 = ~n293 & n303;
  assign n305 = n293 & ~n303;
  assign n306 = ~n304 & ~n305;
  assign n307 = ~n292 & n306;
  assign n308 = n292 & ~n306;
  assign n309 = ~n307 & ~n308;
  assign n310 = ~n291 & ~n309;
  assign n311 = n291 & n309;
  assign n312 = ~n310 & ~n311;
  assign n313 = ~n220 & ~n225;
  assign n314 = n312 & ~n313;
  assign n315 = ~n312 & n313;
  assign n316 = ~n314 & ~n315;
  assign n317 = ~n264 & n316;
  assign n318 = n264 & ~n316;
  assign n319 = ~n317 & ~n318;
  assign n320 = ~n263 & n319;
  assign n321 = ~n314 & ~n317;
  assign n322 = ~n307 & ~n311;
  assign n323 = ~n287 & ~n289;
  assign n324 = ~n269 & ~n275;
  assign n325 = ~n279 & ~n283;
  assign n326 = n296 & ~n325;
  assign n327 = ~n296 & n325;
  assign n328 = ~n326 & ~n327;
  assign n329 = ~n324 & n328;
  assign n330 = n324 & ~n328;
  assign n331 = ~n329 & ~n330;
  assign n332 = ~n323 & n331;
  assign n333 = n323 & ~n331;
  assign n334 = ~n332 & ~n333;
  assign n335 = ~n301 & ~n304;
  assign n336 = pi03 & pi15;
  assign n337 = n270 & n336;
  assign n338 = pi02 & pi15;
  assign n339 = ~n268 & ~n338;
  assign n340 = ~n337 & ~n339;
  assign n341 = pi04 & pi13;
  assign n342 = ~n340 & ~n341;
  assign n343 = n340 & n341;
  assign n344 = ~n342 & ~n343;
  assign n345 = pi06 & pi12;
  assign n346 = n278 & n345;
  assign n347 = pi05 & pi12;
  assign n348 = pi06 & pi11;
  assign n349 = ~n347 & ~n348;
  assign n350 = ~n346 & ~n349;
  assign n351 = pi07 & pi10;
  assign n352 = n350 & n351;
  assign n353 = ~n350 & ~n351;
  assign n354 = ~n352 & ~n353;
  assign n355 = ~n344 & ~n354;
  assign n356 = n344 & n354;
  assign n357 = ~n355 & ~n356;
  assign n358 = ~n335 & n357;
  assign n359 = n335 & ~n357;
  assign n360 = ~n358 & ~n359;
  assign n361 = n334 & n360;
  assign n362 = ~n334 & ~n360;
  assign n363 = ~n361 & ~n362;
  assign n364 = ~n322 & n363;
  assign n365 = n322 & ~n363;
  assign n366 = ~n364 & ~n365;
  assign n367 = n321 & ~n366;
  assign n368 = ~n321 & n366;
  assign n369 = ~n367 & ~n368;
  assign n370 = n320 & n369;
  assign n371 = ~n364 & ~n368;
  assign n372 = ~n332 & ~n361;
  assign n373 = ~n356 & ~n358;
  assign n374 = ~n337 & ~n343;
  assign n375 = n237 & n348;
  assign n376 = pi07 & pi11;
  assign n377 = ~n345 & ~n376;
  assign n378 = ~n375 & ~n377;
  assign n379 = ~n374 & n378;
  assign n380 = n374 & ~n378;
  assign n381 = ~n379 & ~n380;
  assign n382 = ~n373 & n381;
  assign n383 = n373 & ~n381;
  assign n384 = ~n382 & ~n383;
  assign n385 = ~n326 & ~n329;
  assign n386 = pi04 & pi14;
  assign n387 = n336 & n386;
  assign n388 = ~n336 & ~n386;
  assign n389 = ~n387 & ~n388;
  assign n390 = pi05 & pi13;
  assign n391 = n389 & n390;
  assign n392 = ~n389 & ~n390;
  assign n393 = ~n391 & ~n392;
  assign n394 = ~n346 & ~n352;
  assign n395 = n393 & ~n394;
  assign n396 = ~n393 & n394;
  assign n397 = ~n395 & ~n396;
  assign n398 = ~n385 & n397;
  assign n399 = n385 & ~n397;
  assign n400 = ~n398 & ~n399;
  assign n401 = n384 & n400;
  assign n402 = ~n384 & ~n400;
  assign n403 = ~n401 & ~n402;
  assign n404 = ~n372 & n403;
  assign n405 = n372 & ~n403;
  assign n406 = ~n404 & ~n405;
  assign n407 = ~n371 & n406;
  assign n408 = n371 & ~n406;
  assign n409 = ~n407 & ~n408;
  assign n410 = n370 & n409;
  assign n411 = ~n404 & ~n407;
  assign n412 = ~n382 & ~n401;
  assign n413 = ~n395 & ~n398;
  assign n414 = pi05 & pi15;
  assign n415 = n386 & n414;
  assign n416 = pi04 & pi15;
  assign n417 = pi05 & pi14;
  assign n418 = ~n416 & ~n417;
  assign n419 = ~n415 & ~n418;
  assign n420 = pi06 & pi13;
  assign n421 = n419 & n420;
  assign n422 = ~n419 & ~n420;
  assign n423 = ~n421 & ~n422;
  assign n424 = ~n413 & n423;
  assign n425 = n413 & ~n423;
  assign n426 = ~n424 & ~n425;
  assign n427 = ~n375 & ~n379;
  assign n428 = ~n387 & ~n391;
  assign n429 = n237 & ~n428;
  assign n430 = ~n237 & n428;
  assign n431 = ~n429 & ~n430;
  assign n432 = ~n427 & n431;
  assign n433 = n427 & ~n431;
  assign n434 = ~n432 & ~n433;
  assign n435 = n426 & n434;
  assign n436 = ~n426 & ~n434;
  assign n437 = ~n435 & ~n436;
  assign n438 = ~n412 & n437;
  assign n439 = n412 & ~n437;
  assign n440 = ~n438 & ~n439;
  assign n441 = ~n411 & n440;
  assign n442 = n411 & ~n440;
  assign n443 = ~n441 & ~n442;
  assign n444 = n410 & n443;
  assign n445 = ~n438 & ~n441;
  assign n446 = ~n424 & ~n435;
  assign n447 = ~n429 & ~n432;
  assign n448 = ~n415 & ~n421;
  assign n449 = pi06 & pi14;
  assign n450 = n414 & n449;
  assign n451 = ~n414 & ~n449;
  assign n452 = ~n450 & ~n451;
  assign n453 = pi07 & pi13;
  assign n454 = n452 & n453;
  assign n455 = ~n452 & ~n453;
  assign n456 = ~n454 & ~n455;
  assign n457 = ~n448 & n456;
  assign n458 = n448 & ~n456;
  assign n459 = ~n457 & ~n458;
  assign n460 = ~n447 & n459;
  assign n461 = n447 & ~n459;
  assign n462 = ~n460 & ~n461;
  assign n463 = ~n446 & n462;
  assign n464 = n446 & ~n462;
  assign n465 = ~n463 & ~n464;
  assign n466 = ~n445 & n465;
  assign n467 = n445 & ~n465;
  assign n468 = ~n466 & ~n467;
  assign n469 = n444 & n468;
  assign n470 = ~n463 & ~n466;
  assign n471 = ~n457 & ~n460;
  assign n472 = ~n450 & ~n454;
  assign n473 = pi07 & pi14;
  assign n474 = ~n295 & ~n473;
  assign n475 = n295 & n473;
  assign n476 = ~n474 & ~n475;
  assign n477 = ~n472 & n476;
  assign n478 = n472 & ~n476;
  assign n479 = ~n477 & ~n478;
  assign n480 = ~n471 & n479;
  assign n481 = n471 & ~n479;
  assign n482 = ~n480 & ~n481;
  assign n483 = ~n470 & n482;
  assign n484 = n470 & ~n482;
  assign n485 = ~n483 & ~n484;
  assign n486 = n469 & n485;
  assign n487 = ~n480 & ~n483;
  assign n488 = pi07 & pi15;
  assign n489 = ~n449 & ~n477;
  assign n490 = n488 & ~n489;
  assign n491 = ~n477 & ~n488;
  assign n492 = ~n490 & ~n491;
  assign n493 = ~n487 & n492;
  assign n494 = n487 & ~n492;
  assign n495 = ~n493 & ~n494;
  assign n496 = n486 & n495;
  assign n497 = ~n490 & ~n493;
  assign n498 = ~n496 & n497;
  assign n499 = ~n486 & ~n495;
  assign n500 = ~n496 & ~n499;
  assign n501 = ~n469 & ~n485;
  assign n502 = ~n486 & ~n501;
  assign n503 = ~n444 & ~n468;
  assign n504 = ~n469 & ~n503;
  assign n505 = ~n410 & ~n443;
  assign n506 = ~n444 & ~n505;
  assign n507 = ~n370 & ~n409;
  assign n508 = ~n410 & ~n507;
  assign n509 = ~n320 & ~n369;
  assign n510 = ~n370 & ~n509;
  assign n511 = ~pi23 & ~n258;
  assign n512 = ~n261 & ~n511;
  assign n513 = ~n319 & ~n512;
  assign n514 = ~n320 & ~n513;
  assign n515 = ~n258 & ~n261;
  assign n516 = pi23 & ~n515;
  assign n517 = ~pi23 & n515;
  assign n518 = ~n516 & ~n517;
  assign n519 = ~n203 & ~n204;
  assign n520 = pi22 & ~n519;
  assign n521 = ~n204 & ~n260;
  assign n522 = ~n520 & ~n521;
  assign n523 = ~n199 & ~n200;
  assign n524 = pi21 & ~n523;
  assign n525 = ~pi21 & n523;
  assign n526 = ~n524 & ~n525;
  assign n527 = ~n191 & ~n194;
  assign n528 = pi20 & ~n527;
  assign n529 = ~pi20 & n527;
  assign n530 = ~n528 & ~n529;
  assign n531 = ~n183 & ~n186;
  assign n532 = pi19 & ~n531;
  assign n533 = ~pi19 & n531;
  assign n534 = ~n532 & ~n533;
  assign n535 = ~n175 & ~n178;
  assign n536 = pi18 & ~n535;
  assign n537 = ~n175 & ~n180;
  assign n538 = ~n536 & ~n537;
  assign po00 = ~n498;
  assign po01 = n500;
  assign po02 = n502;
  assign po03 = n504;
  assign po04 = n506;
  assign po05 = n508;
  assign po06 = n510;
  assign po07 = n514;
  assign po08 = ~n518;
  assign po09 = ~n522;
  assign po10 = ~n526;
  assign po11 = ~n530;
  assign po12 = ~n534;
  assign po13 = ~n538;
  assign po14 = 1'b0;
  assign po15 = 1'b0;
endmodule
