module adder_i48_o25 (a,b,r);
input [23:0] a,b;
output [24:0] r;

assign r = a+b;

endmodule

