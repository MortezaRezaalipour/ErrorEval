// Benchmark "circuit" written by ABC on Sat Nov 28 04:42:34 2020

module circuit ( 
    g0, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15,
    g963, g962, g961, g960, g959, g958, g957, g956, g955, g954, g953, g952,
    g951, g950, g949, g948, g947, g946  );
  input  g0, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14,
    g15;
  output g963, g962, g961, g960, g959, g958, g957, g956, g955, g954, g953,
    g952, g951, g950, g949, g948, g947, g946;
  wire g16, g17, g18, g19, g20, g21, g22, g23, g24, g25, g26, g27, g28, g29,
    g30, g31, g32, g33, g34, g35, g36, g37, g38, g39, g40, g41, g42, g43,
    g44, g45, g46, g47, g48, g49, g50, g51, g52, g53, g54, g55, g56, g57,
    g58, g59, g60, g61, g62, g63, g64, g65, g66, g67, g68, g69, g70, g71,
    g72, g73, g74, g75, g76, g77, g78, g79, g80, g81, g82, g83, g84, g85,
    g86, g87, g88, g89, g90, g91, g92, g93, g94, g95, g96, g97, g98, g99,
    g100, g101, g102, g103, g104, g105, g106, g107, g108, g109, g110, g111,
    g112, g113, g114, g115, g116, g117, g118, g119, g120, g121, g122, g123,
    g124, g125, g126, g127, g128, g129, g130, g131, g132, g133, g134, g135,
    g136, g137, g138, g139, g140, g141, g142, g143, g144, g145, g146, g147,
    g148, g149, g150, g151, g152, g153, g154, g155, g156, g157, g158, g159,
    g160, g161, g162, g163, g164, g165, g166, g167, g168, g169, g170, g171,
    g172, g173, g174, g175, g176, g177, g178, g179, g180, g181, g182, g183,
    g184, g185, g186, g187, g188, g189, g190, g191, g192, g193, g194, g195,
    g196, g197, g198, g199, g200, g201, g202, g203, g204, g205, g206, g207,
    g208, g209, g210, g211, g212, g213, g214, g215, g216, g217, g218, g219,
    g220, g221, g222, g223, g224, g225, g226, g227, g228, g229, g230, g231,
    g232, g233, g234, g235, g236, g237, g238, g239, g240, g241, g242, g243,
    g244, g245, g246, g247, g248, g249, g250, g251, g252, g253, g254, g255,
    g256, g257, g258, g259, g260, g261, g262, g263, g264, g265, g266, g267,
    g268, g269, g270, g271, g272, g273, g274, g275, g276, g277, g278, g279,
    g280, g281, g282, g283, g284, g285, g286, g287, g288, g289, g290, g291,
    g292, g293, g294, g295, g296, g297, g298, g299, g300, g301, g302, g303,
    g304, g305, g306, g307, g308, g309, g310, g311, g312, g313, g314, g315,
    g316, g317, g318, g319, g320, g321, g322, g323, g324, g325, g326, g327,
    g328, g329, g330, g331, g332, g333, g334, g335, g336, g337, g338, g339,
    g340, g341, g342, g343, g344, g345, g346, g347, g348, g349, g350, g351,
    g352, g353, g354, g355, g356, g357, g358, g359, g360, g361, g362, g363,
    g364, g365, g366, g367, g368, g369, g370, g371, g372, g373, g374, g375,
    g376, g377, g378, g379, g380, g381, g382, g383, g384, g385, g386, g387,
    g388, g389, g390, g391, g392, g393, g394, g395, g396, g397, g398, g399,
    g400, g401, g402, g403, g404, g405, g406, g407, g408, g409, g410, g411,
    g412, g413, g414, g415, g416, g417, g418, g419, g420, g421, g422, g423,
    g424, g425, g426, g427, g428, g429, g430, g431, g432, g433, g434, g435,
    g436, g437, g438, g439, g440, g441, g442, g443, g444, g445, g446, g447,
    g448, g449, g450, g451, g452, g453, g454, g455, g456, g457, g458, g459,
    g460, g461, g462, g463, g464, g465, g466, g467, g468, g469, g470, g471,
    g472, g473, g474, g475, g476, g477, g478, g479, g480, g481, g482, g483,
    g484, g485, g486, g487, g488, g489, g490, g491, g492, g493, g494, g495,
    g496, g497, g498, g499, g500, g501, g502, g503, g504, g505, g506, g507,
    g508, g509, g510, g511, g512, g513, g514, g515, g516, g517, g518, g519,
    g520, g521, g522, g523, g524, g525, g526, g527, g528, g529, g530, g531,
    g532, g533, g534, g535, g536, g537, g538, g539, g540, g541, g542, g543,
    g544, g545, g546, g547, g548, g549, g550, g551, g552, g553, g554, g555,
    g556, g557, g558, g559, g560, g561, g562, g563, g564, g565, g566, g567,
    g568, g569, g570, g571, g572, g573, g574, g575, g576, g577, g578, g579,
    g580, g581, g582, g583, g584, g585, g586, g587, g588, g589, g590, g591,
    g592, g593, g594, g595, g596, g597, g598, g599, g600, g601, g602, g603,
    g604, g605, g606, g607, g608, g609, g610, g611, g612, g613, g614, g615,
    g616, g617, g618, g619, g620, g621, g622, g623, g624, g625, g626, g627,
    g628, g629, g630, g631, g632, g633, g634, g635, g636, g637, g638, g639,
    g640, g641, g642, g643, g644, g645, g646, g647, g648, g649, g650, g651,
    g652, g653, g654, g655, g656, g657, g658, g659, g660, g661, g662, g663,
    g664, g665, g666, g667, g668, g669, g670, g671, g672, g673, g674, g675,
    g676, g677, g678, g679, g680, g681, g682, g683, g684, g685, g686, g687,
    g688, g689, g690, g691, g692, g693, g694, g695, g696, g697, g698, g699,
    g700, g701, g702, g703, g704, g705, g706, g707, g708, g709, g710, g711,
    g712, g713, g714, g715, g716, g717, g718, g719, g720, g721, g722, g723,
    g724, g725, g726, g727, g728, g729, g730, g731, g732, g733, g734, g735,
    g736, g737, g738, g739, g740, g741, g742, g743, g744, g745, g746, g747,
    g748, g749, g750, g751, g752, g753, g754, g755, g756, g757, g758, g759,
    g760, g761, g762, g763, g764, g765, g766, g767, g768, g769, g770, g771,
    g772, g773, g774, g775, g776, g777, g778, g779, g780, g781, g782, g783,
    g784, g785, g786, g787, g788, g789, g790, g791, g792, g793, g794, g795,
    g796, g797, g798, g799, g800, g801, g802, g803, g804, g805, g806, g807,
    g808, g809, g810, g811, g812, g813, g814, g815, g816, g817, g818, g819,
    g820, g821, g822, g823, g824, g825, g826, g827, g828, g829, g830, g831,
    g832, g833, g834, g835, g836, g837, g838, g839, g840, g841, g842, g843,
    g844, g845, g846, g847, g848, g849, g850, g851, g852, g853, g854, g855,
    g856, g857, g858, g859, g860, g861, g862, g863, g864, g865, g866, g867,
    g868, g869, g870, g871, g872, g873, g874, g875, g876, g877, g878, g879,
    g880, g881, g882, g883, g884, g885, g886, g887, g888, g889, g890, g891,
    g892, g893, g894, g895, g896, g897, g898, g899, g900, g901, g902, g903,
    g904, g905, g906, g907, g908, g909, g910, g911, g912, g913, g914, g915,
    g916, g917, g918, g919, g920, g921, g922, g923, g924, g925, g926, g927,
    g928, g929, g930, g931, g932, g933, g934, g935, g936, g937, g938, g939,
    g940, g941, g942, g943, g944, g945;
  assign g16 = ~g15;
  assign g17 = ~g7 & ~g16;
  assign g18 = ~g17;
  assign g19 = ~g7 | ~g16;
  assign g20 = ~g18 | ~g19;
  assign g21 = ~g14;
  assign g22 = ~g6 | ~g21;
  assign g23 = ~g6;
  assign g24 = ~g14 | ~g23;
  assign g25 = ~g22 | ~g24;
  assign g26 = ~g18 | ~g25;
  assign g27 = ~g25;
  assign g28 = ~g17 | ~g27;
  assign g29 = ~g26 | ~g28;
  assign g30 = ~g13;
  assign g31 = ~g5 | ~g30;
  assign g32 = ~g5;
  assign g33 = ~g13 | ~g32;
  assign g34 = ~g31 | ~g33;
  assign g35 = ~g6 | ~g18;
  assign g36 = ~g17 | ~g23;
  assign g37 = ~g21 | ~g36;
  assign g38 = ~g35 | ~g37;
  assign g39 = ~g34 | ~g38;
  assign g40 = ~g34;
  assign g41 = ~g38;
  assign g42 = ~g40 | ~g41;
  assign g43 = ~g39 | ~g42;
  assign g44 = ~g12;
  assign g45 = ~g4 | ~g44;
  assign g46 = ~g4;
  assign g47 = ~g12 | ~g46;
  assign g48 = ~g45 | ~g47;
  assign g49 = ~g5 | ~g38;
  assign g50 = ~g32 | ~g41;
  assign g51 = ~g30 | ~g50;
  assign g52 = ~g49 | ~g51;
  assign g53 = ~g48 | ~g52;
  assign g54 = ~g48;
  assign g55 = ~g52;
  assign g56 = ~g54 | ~g55;
  assign g57 = ~g53 | ~g56;
  assign g58 = ~g11;
  assign g59 = ~g3 | ~g58;
  assign g60 = ~g3;
  assign g61 = ~g11 | ~g60;
  assign g62 = ~g59 | ~g61;
  assign g63 = ~g4 | ~g52;
  assign g64 = ~g46 | ~g55;
  assign g65 = ~g44 | ~g64;
  assign g66 = ~g63 | ~g65;
  assign g67 = ~g62 | ~g66;
  assign g68 = ~g62;
  assign g69 = ~g66;
  assign g70 = ~g68 | ~g69;
  assign g71 = ~g67 | ~g70;
  assign g72 = ~g10;
  assign g73 = ~g2 | ~g72;
  assign g74 = ~g2;
  assign g75 = ~g10 | ~g74;
  assign g76 = ~g73 | ~g75;
  assign g77 = ~g3 | ~g66;
  assign g78 = ~g60 | ~g69;
  assign g79 = ~g58 | ~g78;
  assign g80 = ~g77 | ~g79;
  assign g81 = ~g76 | ~g80;
  assign g82 = ~g76;
  assign g83 = ~g80;
  assign g84 = ~g82 | ~g83;
  assign g85 = ~g81 | ~g84;
  assign g86 = ~g9;
  assign g87 = ~g1 | ~g86;
  assign g88 = ~g1;
  assign g89 = ~g9 | ~g88;
  assign g90 = ~g87 | ~g89;
  assign g91 = ~g2 | ~g80;
  assign g92 = ~g74 | ~g83;
  assign g93 = ~g72 | ~g92;
  assign g94 = ~g91 | ~g93;
  assign g95 = ~g90 | ~g94;
  assign g96 = ~g90;
  assign g97 = ~g94;
  assign g98 = ~g96 | ~g97;
  assign g99 = ~g95 | ~g98;
  assign g100 = ~g8;
  assign g101 = ~g0 | ~g100;
  assign g102 = ~g0;
  assign g103 = ~g8 | ~g102;
  assign g104 = ~g101 | ~g103;
  assign g105 = ~g1 | ~g94;
  assign g106 = ~g88 | ~g97;
  assign g107 = ~g86 | ~g106;
  assign g108 = ~g105 | ~g107;
  assign g109 = ~g104 | ~g108;
  assign g110 = ~g104;
  assign g111 = ~g108;
  assign g112 = ~g110 | ~g111;
  assign g113 = ~g109 | ~g112;
  assign g114 = ~g0 | ~g108;
  assign g115 = ~g102 | ~g111;
  assign g116 = ~g100 | ~g115;
  assign g117 = ~g114 | ~g116;
  assign g118 = ~g104 | ~g117;
  assign g119 = ~g117;
  assign g120 = ~g110 | ~g119;
  assign g121 = ~g118 | ~g120;
  assign g122 = ~g20 | ~g20;
  assign g123 = ~g43 | ~g121;
  assign g124 = ~g71 | ~g99;
  assign g125 = ~g57 | ~g113;
  assign g126 = ~g71 | ~g85;
  assign g127 = ~g126;
  assign g128 = ~g43 | ~g113;
  assign g129 = ~g127 | ~g128;
  assign g130 = ~g128;
  assign g131 = ~g126 | ~g130;
  assign g132 = ~g129 | ~g131;
  assign g133 = ~g71 | ~g71;
  assign g134 = ~g133;
  assign g135 = ~g29 | ~g113;
  assign g136 = ~g135;
  assign g137 = ~g127 | ~g130;
  assign g138 = ~g20 | ~g121;
  assign g139 = ~g43 | ~g99;
  assign g140 = ~g20 | ~g121;
  assign g141 = ~g20 | ~g113;
  assign g142 = ~g29 | ~g99;
  assign g143 = ~g57 | ~g85;
  assign g144 = ~g43 | ~g99;
  assign g145 = ~g144;
  assign g146 = ~g143 | ~g145;
  assign g147 = ~g57 | ~g85;
  assign g148 = ~g147;
  assign g149 = ~g43 | ~g113;
  assign g150 = ~g71 | ~g85;
  assign g151 = ~g130 | ~g150;
  assign g152 = ~g150;
  assign g153 = ~g149 | ~g152;
  assign g154 = ~g151 | ~g153;
  assign g155 = ~g145 | ~g148;
  assign g156 = ~g99 | ~g155;
  assign g157 = ~g156;
  assign g158 = ~g57 | ~g157;
  assign g159 = ~g154 | ~g158;
  assign g160 = ~g29 | ~g121;
  assign g161 = ~g57 | ~g99;
  assign g162 = ~g161;
  assign g163 = ~g160 | ~g162;
  assign g164 = ~g29 | ~g121;
  assign g165 = ~g164;
  assign g166 = ~g140;
  assign g167 = ~g57 | ~g71;
  assign g168 = ~g167;
  assign g169 = ~g43 | ~g71;
  assign g170 = ~g169;
  assign g171 = ~g43 | ~g71;
  assign g172 = ~g171;
  assign g173 = ~g29 | ~g85;
  assign g174 = ~g172 | ~g173;
  assign g175 = ~g173;
  assign g176 = ~g171 | ~g175;
  assign g177 = ~g174 | ~g176;
  assign g178 = ~g170 | ~g177;
  assign g179 = ~g172 | ~g175;
  assign g180 = ~g178 | ~g179;
  assign g181 = ~g57 | ~g113;
  assign g182 = ~g181;
  assign g183 = ~g71 | ~g99;
  assign g184 = ~g182 | ~g183;
  assign g185 = ~g183;
  assign g186 = ~g181 | ~g185;
  assign g187 = ~g184 | ~g186;
  assign g188 = ~g149 | ~g150;
  assign g189 = ~g188;
  assign g190 = ~g85 | ~g85;
  assign g191 = ~g189 | ~g190;
  assign g192 = ~g190;
  assign g193 = ~g188 | ~g192;
  assign g194 = ~g191 | ~g193;
  assign g195 = ~g43 | ~g121;
  assign g196 = ~g194 | ~g195;
  assign g197 = ~g195;
  assign g198 = ~g194;
  assign g199 = ~g197 | ~g198;
  assign g200 = ~g196 | ~g199;
  assign g201 = ~g200;
  assign g202 = ~g29 | ~g85;
  assign g203 = ~g202;
  assign g204 = ~g20 | ~g99;
  assign g205 = ~g204;
  assign g206 = ~g203 | ~g205;
  assign g207 = ~g206;
  assign g208 = ~g20 | ~g113;
  assign g209 = ~g208;
  assign g210 = ~g43 | ~g85;
  assign g211 = ~g210;
  assign g212 = ~g43 | ~g85;
  assign g213 = ~g29 | ~g99;
  assign g214 = ~g211 | ~g213;
  assign g215 = ~g213;
  assign g216 = ~g212 | ~g215;
  assign g217 = ~g214 | ~g216;
  assign g218 = ~g211 | ~g217;
  assign g219 = ~g211 | ~g215;
  assign g220 = ~g218 | ~g219;
  assign g221 = ~g220;
  assign g222 = ~g210 | ~g217;
  assign g223 = ~g217;
  assign g224 = ~g211 | ~g223;
  assign g225 = ~g222 | ~g224;
  assign g226 = ~g225;
  assign g227 = ~g169 | ~g177;
  assign g228 = ~g177;
  assign g229 = ~g170 | ~g228;
  assign g230 = ~g227 | ~g229;
  assign g231 = ~g43 | ~g57;
  assign g232 = ~g231;
  assign g233 = ~g29 | ~g71;
  assign g234 = ~g43 | ~g57;
  assign g235 = ~g232 | ~g233;
  assign g236 = ~g57 | ~g57;
  assign g237 = ~g236;
  assign g238 = ~g20 | ~g85;
  assign g239 = ~g29 | ~g71;
  assign g240 = ~g239;
  assign g241 = ~g203 | ~g204;
  assign g242 = ~g202 | ~g205;
  assign g243 = ~g241 | ~g242;
  assign g244 = ~g20 | ~g99;
  assign g245 = ~g243 | ~g244;
  assign g246 = ~g243;
  assign g247 = ~g244;
  assign g248 = ~g246 | ~g247;
  assign g249 = ~g245 | ~g248;
  assign g250 = ~g243 | ~g247;
  assign g251 = ~g230;
  assign g252 = ~g29 | ~g57;
  assign g253 = ~g20 | ~g71;
  assign g254 = ~g253;
  assign g255 = ~g238 | ~g240;
  assign g256 = ~g20 | ~g85;
  assign g257 = ~g256;
  assign g258 = ~g249;
  assign g259 = ~g43 | ~g43;
  assign g260 = ~g259;
  assign g261 = ~g29 | ~g57;
  assign g262 = ~g260 | ~g261;
  assign g263 = ~g261;
  assign g264 = ~g259 | ~g263;
  assign g265 = ~g262 | ~g264;
  assign g266 = ~g29 | ~g29;
  assign g267 = ~g266;
  assign g268 = ~g20 | ~g43;
  assign g269 = ~g20 | ~g57;
  assign g270 = ~g29 | ~g43;
  assign g271 = ~g270;
  assign g272 = ~g260 | ~g263;
  assign g273 = ~g20 | ~g57;
  assign g274 = ~g273;
  assign g275 = ~g29 | ~g43;
  assign g276 = ~g271 | ~g274;
  assign g277 = ~g276;
  assign g278 = ~g252 | ~g254;
  assign g279 = ~g253 | ~g263;
  assign g280 = ~g278 | ~g279;
  assign g281 = ~g20 | ~g71;
  assign g282 = ~g280 | ~g281;
  assign g283 = ~g280;
  assign g284 = ~g254 | ~g283;
  assign g285 = ~g282 | ~g284;
  assign g286 = ~g277 | ~g285;
  assign g287 = ~g254 | ~g280;
  assign g288 = ~g286 | ~g287;
  assign g289 = ~g288;
  assign g290 = ~g276 | ~g285;
  assign g291 = ~g285;
  assign g292 = ~g277 | ~g291;
  assign g293 = ~g290 | ~g292;
  assign g294 = ~g293;
  assign g295 = ~g269 | ~g271;
  assign g296 = ~g270 | ~g274;
  assign g297 = ~g295 | ~g296;
  assign g298 = ~g271 | ~g273;
  assign g299 = ~g274 | ~g275;
  assign g300 = ~g298 | ~g299;
  assign g301 = ~g300;
  assign g302 = ~g20 | ~g29;
  assign g303 = ~g302;
  assign g304 = ~g303 | ~g303;
  assign g305 = ~g304;
  assign g306 = ~g267 | ~g268;
  assign g307 = ~g20 | ~g43;
  assign g308 = ~g307;
  assign g309 = ~g85 | ~g99;
  assign g310 = ~g309;
  assign g311 = ~g71 | ~g113;
  assign g312 = ~g310 | ~g311;
  assign g313 = ~g71 | ~g113;
  assign g314 = ~g313;
  assign g315 = ~g182 | ~g185;
  assign g316 = ~g57 | ~g121;
  assign g317 = ~g85 | ~g99;
  assign g318 = ~g310 | ~g316;
  assign g319 = ~g57 | ~g121;
  assign g320 = ~g319;
  assign g321 = ~g195 | ~g198;
  assign g322 = ~g193 | ~g321;
  assign g323 = ~g322;
  assign g324 = ~g85 | ~g113;
  assign g325 = ~g324;
  assign g326 = ~g310 | ~g314;
  assign g327 = ~g71 | ~g121;
  assign g328 = ~g99 | ~g99;
  assign g329 = ~g328;
  assign g330 = ~g327 | ~g329;
  assign g331 = ~g71 | ~g121;
  assign g332 = ~g331;
  assign g333 = ~g99 | ~g113;
  assign g334 = ~g85 | ~g121;
  assign g335 = ~g99 | ~g113;
  assign g336 = ~g335;
  assign g337 = ~g334 | ~g336;
  assign g338 = ~g85 | ~g121;
  assign g339 = ~g338;
  assign g340 = ~g99 | ~g121;
  assign g341 = ~g113 | ~g113;
  assign g342 = ~g341;
  assign g343 = ~g340 | ~g342;
  assign g344 = ~g99 | ~g121;
  assign g345 = ~g344;
  assign g346 = ~g113 | ~g121;
  assign g347 = ~g113 | ~g121;
  assign g348 = ~g347;
  assign g349 = ~g346 | ~g347;
  assign g350 = ~g121 | ~g121;
  assign g351 = ~g350;
  assign g352 = ~g347 & ~g348;
  assign g353 = ~g154 & ~g158;
  assign g354 = ~g167 & ~g168;
  assign g355 = ~g324 & ~g325;
  assign g356 = ~g135 & ~g136;
  assign g357 = ~g124 | ~g197;
  assign g358 = ~g123 | ~g185;
  assign g359 = ~g357 | ~g358;
  assign g360 = ~g125 | ~g359;
  assign g361 = ~g359;
  assign g362 = ~g182 | ~g361;
  assign g363 = ~g360 | ~g362;
  assign g364 = ~g134 | ~g356;
  assign g365 = ~g363;
  assign g366 = ~g139 | ~g166;
  assign g367 = ~g138 | ~g145;
  assign g368 = ~g366 | ~g367;
  assign g369 = ~g368;
  assign g370 = ~g140 | ~g369;
  assign g371 = ~g367 | ~g370;
  assign g372 = ~g371;
  assign g373 = ~g209 | ~g215;
  assign g374 = ~g373;
  assign g375 = ~g144 | ~g148;
  assign g376 = ~g146 | ~g375;
  assign g377 = ~g147 | ~g376;
  assign g378 = ~g376;
  assign g379 = ~g148 | ~g378;
  assign g380 = ~g377 | ~g379;
  assign g381 = ~g374 | ~g380;
  assign g382 = ~g148 | ~g376;
  assign g383 = ~g381 | ~g382;
  assign g384 = ~g161 | ~g165;
  assign g385 = ~g163 | ~g384;
  assign g386 = ~g164 | ~g385;
  assign g387 = ~g385;
  assign g388 = ~g165 | ~g387;
  assign g389 = ~g386 | ~g388;
  assign g390 = ~g389;
  assign g391 = ~g140 | ~g368;
  assign g392 = ~g166 | ~g369;
  assign g393 = ~g391 | ~g392;
  assign g394 = ~g133 | ~g356;
  assign g395 = ~g356;
  assign g396 = ~g134 | ~g395;
  assign g397 = ~g394 | ~g396;
  assign g398 = ~g397;
  assign g399 = ~g393 | ~g398;
  assign g400 = ~g393;
  assign g401 = ~g397 | ~g400;
  assign g402 = ~g399 | ~g401;
  assign g403 = ~g180 | ~g354;
  assign g404 = ~g393 | ~g397;
  assign g405 = ~g164 | ~g387;
  assign g406 = ~g163 | ~g405;
  assign g407 = ~g187 | ~g406;
  assign g408 = ~g187 & ~g406;
  assign g409 = ~g408;
  assign g410 = ~g407 | ~g409;
  assign g411 = ~g410;
  assign g412 = ~g142 | ~g209;
  assign g413 = ~g141 | ~g215;
  assign g414 = ~g412 | ~g413;
  assign g415 = ~g208 | ~g414;
  assign g416 = ~g414;
  assign g417 = ~g209 | ~g416;
  assign g418 = ~g415 | ~g417;
  assign g419 = ~g207 | ~g418;
  assign g420 = ~g209 | ~g414;
  assign g421 = ~g419 | ~g420;
  assign g422 = ~g421;
  assign g423 = ~g220 | ~g422;
  assign g424 = ~g221 | ~g421;
  assign g425 = ~g423 | ~g424;
  assign g426 = ~g373 | ~g380;
  assign g427 = ~g380;
  assign g428 = ~g374 | ~g427;
  assign g429 = ~g426 | ~g428;
  assign g430 = ~g425 | ~g429;
  assign g431 = ~g220 | ~g421;
  assign g432 = ~g430 | ~g431;
  assign g433 = ~g429;
  assign g434 = ~g425 | ~g433;
  assign g435 = ~g425;
  assign g436 = ~g429 | ~g435;
  assign g437 = ~g434 | ~g436;
  assign g438 = ~g437;
  assign g439 = ~g206 | ~g418;
  assign g440 = ~g418;
  assign g441 = ~g207 | ~g440;
  assign g442 = ~g439 | ~g441;
  assign g443 = ~g226 | ~g442;
  assign g444 = ~g442;
  assign g445 = ~g225 | ~g444;
  assign g446 = ~g443 | ~g445;
  assign g447 = ~g234 | ~g240;
  assign g448 = ~g235 | ~g447;
  assign g449 = ~g232 | ~g448;
  assign g450 = ~g232 | ~g240;
  assign g451 = ~g449 | ~g450;
  assign g452 = ~g451;
  assign g453 = ~g236 | ~g452;
  assign g454 = ~g237 | ~g451;
  assign g455 = ~g453 | ~g454;
  assign g456 = ~g455;
  assign g457 = ~g230 | ~g456;
  assign g458 = ~g454 | ~g457;
  assign g459 = ~g446 | ~g458;
  assign g460 = ~g225 | ~g442;
  assign g461 = ~g459 | ~g460;
  assign g462 = ~g461;
  assign g463 = ~g180 & ~g354;
  assign g464 = ~g463;
  assign g465 = ~g403 | ~g464;
  assign g466 = ~g240 | ~g257;
  assign g467 = ~g466;
  assign g468 = ~g249 | ~g467;
  assign g469 = ~g250 | ~g468;
  assign g470 = ~g465 | ~g469;
  assign g471 = ~g469;
  assign g472 = ~g465;
  assign g473 = ~g471 | ~g472;
  assign g474 = ~g470 | ~g473;
  assign g475 = ~g446 & ~g458;
  assign g476 = ~g475;
  assign g477 = ~g459 | ~g476;
  assign g478 = ~g477;
  assign g479 = ~g474 | ~g478;
  assign g480 = ~g469 | ~g472;
  assign g481 = ~g479 | ~g480;
  assign g482 = ~g474;
  assign g483 = ~g477 | ~g482;
  assign g484 = ~g479 | ~g483;
  assign g485 = ~g251 | ~g455;
  assign g486 = ~g457 | ~g485;
  assign g487 = ~g254 | ~g263;
  assign g488 = ~g487;
  assign g489 = ~g239 | ~g257;
  assign g490 = ~g255 | ~g489;
  assign g491 = ~g256 | ~g490;
  assign g492 = ~g490;
  assign g493 = ~g257 | ~g492;
  assign g494 = ~g491 | ~g493;
  assign g495 = ~g488 | ~g494;
  assign g496 = ~g257 | ~g490;
  assign g497 = ~g495 | ~g496;
  assign g498 = ~g486 | ~g497;
  assign g499 = ~g497;
  assign g500 = ~g486;
  assign g501 = ~g499 | ~g500;
  assign g502 = ~g498 | ~g501;
  assign g503 = ~g249 | ~g466;
  assign g504 = ~g258 | ~g467;
  assign g505 = ~g503 | ~g504;
  assign g506 = ~g502 | ~g505;
  assign g507 = ~g497 | ~g500;
  assign g508 = ~g506 | ~g507;
  assign g509 = ~g484 | ~g508;
  assign g510 = ~g508;
  assign g511 = ~g484;
  assign g512 = ~g510 | ~g511;
  assign g513 = ~g509 | ~g512;
  assign g514 = ~g505;
  assign g515 = ~g502 | ~g514;
  assign g516 = ~g502;
  assign g517 = ~g505 | ~g516;
  assign g518 = ~g515 | ~g517;
  assign g519 = ~g231 | ~g448;
  assign g520 = ~g448;
  assign g521 = ~g232 | ~g520;
  assign g522 = ~g519 | ~g521;
  assign g523 = ~g267 | ~g308;
  assign g524 = ~g271 | ~g274;
  assign g525 = ~g523 | ~g524;
  assign g526 = ~g265 | ~g525;
  assign g527 = ~g272 | ~g526;
  assign g528 = ~g522 | ~g527;
  assign g529 = ~g522 & ~g527;
  assign g530 = ~g529;
  assign g531 = ~g528 | ~g530;
  assign g532 = ~g531;
  assign g533 = ~g288 | ~g532;
  assign g534 = ~g528 | ~g533;
  assign g535 = ~g518 | ~g534;
  assign g536 = ~g518 & ~g534;
  assign g537 = ~g536;
  assign g538 = ~g535 | ~g537;
  assign g539 = ~g538;
  assign g540 = ~g288 | ~g531;
  assign g541 = ~g289 | ~g532;
  assign g542 = ~g540 | ~g541;
  assign g543 = ~g487 | ~g494;
  assign g544 = ~g494;
  assign g545 = ~g488 | ~g544;
  assign g546 = ~g543 | ~g545;
  assign g547 = ~g546;
  assign g548 = ~g542 | ~g547;
  assign g549 = ~g542;
  assign g550 = ~g546 | ~g549;
  assign g551 = ~g548 | ~g550;
  assign g552 = ~g265 & ~g525;
  assign g553 = ~g552;
  assign g554 = ~g526 | ~g553;
  assign g555 = ~g294 | ~g554;
  assign g556 = ~g554;
  assign g557 = ~g293 | ~g556;
  assign g558 = ~g555 | ~g557;
  assign g559 = ~g558;
  assign g560 = ~g297 | ~g523;
  assign g561 = ~g297 & ~g523;
  assign g562 = ~g561;
  assign g563 = ~g560 | ~g562;
  assign g564 = ~g301 | ~g563;
  assign g565 = ~g563;
  assign g566 = ~g300 | ~g565;
  assign g567 = ~g564 | ~g566;
  assign g568 = ~g266 | ~g308;
  assign g569 = ~g306 | ~g568;
  assign g570 = ~g307 | ~g569;
  assign g571 = ~g569;
  assign g572 = ~g308 | ~g571;
  assign g573 = ~g570 | ~g572;
  assign g574 = ~g305 | ~g573;
  assign g575 = ~g308 | ~g569;
  assign g576 = ~g574 | ~g575;
  assign g577 = ~g567 | ~g576;
  assign g578 = ~g300 | ~g563;
  assign g579 = ~g577 | ~g578;
  assign g580 = ~g559 | ~g579;
  assign g581 = ~g557 | ~g580;
  assign g582 = ~g551 | ~g581;
  assign g583 = ~g542 | ~g546;
  assign g584 = ~g582 | ~g583;
  assign g585 = ~g539 | ~g584;
  assign g586 = ~g535 | ~g585;
  assign g587 = ~g513 | ~g586;
  assign g588 = ~g508 | ~g511;
  assign g589 = ~g587 | ~g588;
  assign g590 = ~g309 | ~g314;
  assign g591 = ~g312 | ~g590;
  assign g592 = ~g313 | ~g591;
  assign g593 = ~g591;
  assign g594 = ~g314 | ~g593;
  assign g595 = ~g592 | ~g594;
  assign g596 = ~g315 | ~g407;
  assign g597 = ~g595 | ~g596;
  assign g598 = ~g595 & ~g596;
  assign g599 = ~g598;
  assign g600 = ~g597 | ~g599;
  assign g601 = ~g317 | ~g320;
  assign g602 = ~g318 | ~g601;
  assign g603 = ~g319 | ~g602;
  assign g604 = ~g602;
  assign g605 = ~g320 | ~g604;
  assign g606 = ~g603 | ~g605;
  assign g607 = ~g606;
  assign g608 = ~g600 | ~g607;
  assign g609 = ~g600;
  assign g610 = ~g606 | ~g609;
  assign g611 = ~g608 | ~g610;
  assign g612 = ~g358 | ~g362;
  assign g613 = ~g323 | ~g612;
  assign g614 = ~g612;
  assign g615 = ~g322 | ~g614;
  assign g616 = ~g613 | ~g615;
  assign g617 = ~g611;
  assign g618 = ~g322 | ~g612;
  assign g619 = ~g597 | ~g610;
  assign g620 = ~g619;
  assign g621 = ~g314 | ~g591;
  assign g622 = ~g326 | ~g621;
  assign g623 = ~g355 | ~g622;
  assign g624 = ~g355 & ~g622;
  assign g625 = ~g624;
  assign g626 = ~g623 | ~g625;
  assign g627 = ~g319 | ~g604;
  assign g628 = ~g318 | ~g627;
  assign g629 = ~g626 | ~g628;
  assign g630 = ~g628;
  assign g631 = ~g626;
  assign g632 = ~g630 | ~g631;
  assign g633 = ~g629 | ~g632;
  assign g634 = ~g328 | ~g332;
  assign g635 = ~g330 | ~g634;
  assign g636 = ~g331 | ~g635;
  assign g637 = ~g635;
  assign g638 = ~g332 | ~g637;
  assign g639 = ~g636 | ~g638;
  assign g640 = ~g639;
  assign g641 = ~g633 | ~g640;
  assign g642 = ~g633;
  assign g643 = ~g639 | ~g642;
  assign g644 = ~g641 | ~g643;
  assign g645 = ~g644;
  assign g646 = ~g331 | ~g637;
  assign g647 = ~g330 | ~g646;
  assign g648 = ~g647;
  assign g649 = ~g333 | ~g648;
  assign g650 = ~g336 | ~g647;
  assign g651 = ~g649 | ~g650;
  assign g652 = ~g651;
  assign g653 = ~g335 | ~g339;
  assign g654 = ~g337 | ~g653;
  assign g655 = ~g338 | ~g654;
  assign g656 = ~g654;
  assign g657 = ~g339 | ~g656;
  assign g658 = ~g655 | ~g657;
  assign g659 = ~g658;
  assign g660 = ~g633 | ~g639;
  assign g661 = ~g628 | ~g631;
  assign g662 = ~g660 | ~g661;
  assign g663 = ~g341 | ~g345;
  assign g664 = ~g343 | ~g663;
  assign g665 = ~g344 | ~g664;
  assign g666 = ~g664;
  assign g667 = ~g345 | ~g666;
  assign g668 = ~g665 | ~g667;
  assign g669 = ~g338 | ~g656;
  assign g670 = ~g337 | ~g669;
  assign g671 = ~g668 | ~g670;
  assign g672 = ~g668 & ~g670;
  assign g673 = ~g672;
  assign g674 = ~g671 | ~g673;
  assign g675 = ~g674;
  assign g676 = ~g344 | ~g666;
  assign g677 = ~g343 | ~g676;
  assign g678 = ~g352 | ~g677;
  assign g679 = ~g352 & ~g677;
  assign g680 = ~g679;
  assign g681 = ~g678 | ~g680;
  assign g682 = ~g681;
  assign g683 = ~g349 | ~g678;
  assign g684 = ~g683;
  assign g685 = ~g350 | ~g684;
  assign g686 = ~g351 | ~g683;
  assign g687 = ~g685 | ~g686;
  assign g688 = ~g687;
  assign g689 = ~g304 | ~g573;
  assign g690 = ~g573;
  assign g691 = ~g305 | ~g690;
  assign g692 = ~g577;
  assign g693 = ~g567 & ~g576;
  assign g694 = ~g558 | ~g579;
  assign g695 = ~g579;
  assign g696 = ~g559 | ~g695;
  assign g697 = ~g582;
  assign g698 = ~g551 & ~g581;
  assign g699 = ~g538 | ~g584;
  assign g700 = ~g584;
  assign g701 = ~g539 | ~g700;
  assign g702 = ~g587;
  assign g703 = ~g513 & ~g586;
  assign g704 = ~g589;
  assign g705 = ~g324 | ~g623;
  assign g706 = ~g167 | ~g403;
  assign g707 = ~g353;
  assign g708 = ~g135 | ~g364;
  assign g709 = ~g132 | ~g708;
  assign g710 = ~g137 | ~g709;
  assign g711 = ~g363 | ~g710;
  assign g712 = ~g710;
  assign g713 = ~g365 | ~g712;
  assign g714 = ~g711 | ~g713;
  assign g715 = ~g132 & ~g708;
  assign g716 = ~g715;
  assign g717 = ~g709 | ~g716;
  assign g718 = ~g371 | ~g717;
  assign g719 = ~g717;
  assign g720 = ~g372 | ~g719;
  assign g721 = ~g718 | ~g720;
  assign g722 = ~g383 | ~g721;
  assign g723 = ~g371 | ~g719;
  assign g724 = ~g722 | ~g723;
  assign g725 = ~g714 | ~g724;
  assign g726 = ~g714 & ~g724;
  assign g727 = ~g726;
  assign g728 = ~g725 | ~g727;
  assign g729 = ~g159 | ~g707;
  assign g730 = ~g390 | ~g729;
  assign g731 = ~g729;
  assign g732 = ~g389 | ~g731;
  assign g733 = ~g730 | ~g732;
  assign g734 = ~g733;
  assign g735 = ~g402 | ~g706;
  assign g736 = ~g404 | ~g735;
  assign g737 = ~g734 | ~g736;
  assign g738 = ~g732 | ~g737;
  assign g739 = ~g728 | ~g738;
  assign g740 = ~g738;
  assign g741 = ~g728;
  assign g742 = ~g740 | ~g741;
  assign g743 = ~g739 | ~g742;
  assign g744 = ~g155 | ~g707;
  assign g745 = ~g410 | ~g744;
  assign g746 = ~g744;
  assign g747 = ~g411 | ~g746;
  assign g748 = ~g745 | ~g747;
  assign g749 = ~g201 | ~g748;
  assign g750 = ~g748;
  assign g751 = ~g200 | ~g750;
  assign g752 = ~g749 | ~g751;
  assign g753 = ~g752;
  assign g754 = ~g743 | ~g753;
  assign g755 = ~g743;
  assign g756 = ~g752 | ~g755;
  assign g757 = ~g754 | ~g756;
  assign g758 = ~g383 & ~g721;
  assign g759 = ~g758;
  assign g760 = ~g722 | ~g759;
  assign g761 = ~g760;
  assign g762 = ~g733 | ~g736;
  assign g763 = ~g736;
  assign g764 = ~g734 | ~g763;
  assign g765 = ~g762 | ~g764;
  assign g766 = ~g432 | ~g765;
  assign g767 = ~g432 & ~g765;
  assign g768 = ~g767;
  assign g769 = ~g766 | ~g768;
  assign g770 = ~g769;
  assign g771 = ~g761 | ~g770;
  assign g772 = ~g766 | ~g771;
  assign g773 = ~g757 | ~g772;
  assign g774 = ~g757 & ~g772;
  assign g775 = ~g774;
  assign g776 = ~g773 | ~g775;
  assign g777 = ~g761 | ~g769;
  assign g778 = ~g760 | ~g770;
  assign g779 = ~g777 | ~g778;
  assign g780 = ~g402 & ~g706;
  assign g781 = ~g780;
  assign g782 = ~g735 | ~g781;
  assign g783 = ~g438 | ~g782;
  assign g784 = ~g782;
  assign g785 = ~g437 | ~g784;
  assign g786 = ~g783 | ~g785;
  assign g787 = ~g786;
  assign g788 = ~g461 | ~g787;
  assign g789 = ~g785 | ~g788;
  assign g790 = ~g779 | ~g789;
  assign g791 = ~g779 & ~g789;
  assign g792 = ~g791;
  assign g793 = ~g790 | ~g792;
  assign g794 = ~g793;
  assign g795 = ~g461 | ~g786;
  assign g796 = ~g462 | ~g787;
  assign g797 = ~g795 | ~g796;
  assign g798 = ~g481 | ~g797;
  assign g799 = ~g481 & ~g797;
  assign g800 = ~g799;
  assign g801 = ~g798 | ~g800;
  assign g802 = ~g801;
  assign g803 = ~g589 | ~g802;
  assign g804 = ~g798 | ~g803;
  assign g805 = ~g794 | ~g804;
  assign g806 = ~g790 | ~g805;
  assign g807 = ~g776 | ~g806;
  assign g808 = ~g806;
  assign g809 = ~g776;
  assign g810 = ~g808 | ~g809;
  assign g811 = ~g200 | ~g748;
  assign g812 = ~g411 | ~g744;
  assign g813 = ~g811 | ~g812;
  assign g814 = ~g616 | ~g813;
  assign g815 = ~g616 & ~g813;
  assign g816 = ~g815;
  assign g817 = ~g814 | ~g816;
  assign g818 = ~g817;
  assign g819 = ~g611 | ~g818;
  assign g820 = ~g617 | ~g817;
  assign g821 = ~g819 | ~g820;
  assign g822 = ~g365 | ~g710;
  assign g823 = ~g725 | ~g822;
  assign g824 = ~g821 | ~g823;
  assign g825 = ~g821 & ~g823;
  assign g826 = ~g825;
  assign g827 = ~g824 | ~g826;
  assign g828 = ~g743 | ~g752;
  assign g829 = ~g738 | ~g741;
  assign g830 = ~g828 | ~g829;
  assign g831 = ~g827 | ~g830;
  assign g832 = ~g830;
  assign g833 = ~g827;
  assign g834 = ~g832 | ~g833;
  assign g835 = ~g831 | ~g834;
  assign g836 = ~g806 | ~g809;
  assign g837 = ~g773 | ~g836;
  assign g838 = ~g835 | ~g837;
  assign g839 = ~g838;
  assign g840 = ~g835 & ~g837;
  assign g841 = ~g618 | ~g814;
  assign g842 = ~g841;
  assign g843 = ~g619 | ~g842;
  assign g844 = ~g620 | ~g841;
  assign g845 = ~g843 | ~g844;
  assign g846 = ~g645 | ~g845;
  assign g847 = ~g845;
  assign g848 = ~g644 | ~g847;
  assign g849 = ~g846 | ~g848;
  assign g850 = ~g617 | ~g818;
  assign g851 = ~g824 | ~g850;
  assign g852 = ~g849 | ~g851;
  assign g853 = ~g849 & ~g851;
  assign g854 = ~g853;
  assign g855 = ~g852 | ~g854;
  assign g856 = ~g830 | ~g833;
  assign g857 = ~g838 | ~g856;
  assign g858 = ~g855 | ~g857;
  assign g859 = ~g857;
  assign g860 = ~g855;
  assign g861 = ~g859 | ~g860;
  assign g862 = ~g651 | ~g705;
  assign g863 = ~g705;
  assign g864 = ~g652 | ~g863;
  assign g865 = ~g862 | ~g864;
  assign g866 = ~g659 | ~g865;
  assign g867 = ~g865;
  assign g868 = ~g658 | ~g867;
  assign g869 = ~g866 | ~g868;
  assign g870 = ~g662 | ~g869;
  assign g871 = ~g662 & ~g869;
  assign g872 = ~g871;
  assign g873 = ~g870 | ~g872;
  assign g874 = ~g644 | ~g845;
  assign g875 = ~g619 | ~g841;
  assign g876 = ~g874 | ~g875;
  assign g877 = ~g873 | ~g876;
  assign g878 = ~g876;
  assign g879 = ~g873;
  assign g880 = ~g878 | ~g879;
  assign g881 = ~g877 | ~g880;
  assign g882 = ~g857 | ~g860;
  assign g883 = ~g852 | ~g882;
  assign g884 = ~g881 | ~g883;
  assign g885 = ~g884;
  assign g886 = ~g881 & ~g883;
  assign g887 = ~g652 | ~g705;
  assign g888 = ~g650 | ~g887;
  assign g889 = ~g674 | ~g888;
  assign g890 = ~g888;
  assign g891 = ~g675 | ~g890;
  assign g892 = ~g889 | ~g891;
  assign g893 = ~g658 | ~g865;
  assign g894 = ~g870 | ~g893;
  assign g895 = ~g892 | ~g894;
  assign g896 = ~g892 & ~g894;
  assign g897 = ~g896;
  assign g898 = ~g895 | ~g897;
  assign g899 = ~g876 | ~g879;
  assign g900 = ~g884 | ~g899;
  assign g901 = ~g898 | ~g900;
  assign g902 = ~g900;
  assign g903 = ~g898;
  assign g904 = ~g902 | ~g903;
  assign g905 = ~g675 | ~g888;
  assign g906 = ~g671 | ~g905;
  assign g907 = ~g681 | ~g906;
  assign g908 = ~g906;
  assign g909 = ~g682 | ~g908;
  assign g910 = ~g907 | ~g909;
  assign g911 = ~g900 | ~g903;
  assign g912 = ~g895 | ~g911;
  assign g913 = ~g910 | ~g912;
  assign g914 = ~g913;
  assign g915 = ~g910 & ~g912;
  assign g916 = ~g682 | ~g906;
  assign g917 = ~g913 | ~g916;
  assign g918 = ~g687 | ~g917;
  assign g919 = ~g917;
  assign g920 = ~g688 | ~g919;
  assign g921 = ~g688 | ~g917;
  assign g922 = ~g686 | ~g921;
  assign g923 = ~g589 | ~g801;
  assign g924 = ~g704 | ~g802;
  assign g925 = ~g793 | ~g804;
  assign g926 = ~g804;
  assign g927 = ~g794 | ~g926;
  assign g928 = ~g122;
  assign g929 = ~g302 & ~g303;
  assign g930 = ~g689 | ~g691;
  assign g931 = ~g692 & ~g693;
  assign g932 = ~g694 | ~g696;
  assign g933 = ~g697 & ~g698;
  assign g934 = ~g699 | ~g701;
  assign g935 = ~g702 & ~g703;
  assign g936 = ~g923 | ~g924;
  assign g937 = ~g925 | ~g927;
  assign g938 = ~g807 | ~g810;
  assign g939 = ~g839 & ~g840;
  assign g940 = ~g858 | ~g861;
  assign g941 = ~g885 & ~g886;
  assign g942 = ~g901 | ~g904;
  assign g943 = ~g914 & ~g915;
  assign g944 = ~g918 | ~g920;
  assign g945 = ~g922;
  assign g946 = g928;
  assign g947 = g929;
  assign g948 = g930;
  assign g949 = g931;
  assign g950 = g932;
  assign g951 = g933;
  assign g952 = g934;
  assign g953 = g935;
  assign g954 = g936;
  assign g955 = g937;
  assign g956 = g938;
  assign g957 = g939;
  assign g958 = g940;
  assign g959 = g941;
  assign g960 = g942;
  assign g961 = g943;
  assign g962 = g944;
  assign g963 = g945;
endmodule


