module adder_i28_o15 (a,b,r);
input [13:0] a,b;
output [14:0] r;

assign r = a+b;

endmodule

