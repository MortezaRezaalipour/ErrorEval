module top(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, po0, po1, po2);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09;
  output po0, po1, po2;
  wire n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82;
  assign n11 = pi00 & ~pi06;
  assign n12 = ~pi00 & pi06;
  assign n13 = ~n11 & ~n12;
  assign n14 = pi02 & ~pi04;
  assign n15 = ~pi02 & pi04;
  assign n16 = ~n14 & ~n15;
  assign n17 = ~n13 & ~n16;
  assign n18 = ~pi02 & ~pi04;
  assign n19 = pi02 & pi04;
  assign n20 = ~n18 & ~n19;
  assign n21 = n13 & ~n20;
  assign n22 = ~n17 & ~n21;
  assign n23 = ~pi00 & pi08;
  assign n24 = pi00 & ~pi08;
  assign n25 = ~n23 & ~n24;
  assign n26 = n22 & ~n25;
  assign n27 = ~n22 & n25;
  assign n28 = ~n26 & ~n27;
  assign n29 = ~pi00 & pi04;
  assign n30 = pi02 & n29;
  assign n31 = pi00 & ~pi04;
  assign n32 = ~pi02 & n31;
  assign n33 = ~n30 & ~n32;
  assign n34 = ~n17 & n33;
  assign n35 = pi00 & ~pi02;
  assign n36 = ~pi01 & pi03;
  assign n37 = ~n35 & n36;
  assign n38 = ~pi00 & pi02;
  assign n39 = pi01 & ~pi03;
  assign n40 = ~n38 & n39;
  assign n41 = ~n37 & ~n40;
  assign n42 = ~pi01 & pi05;
  assign n43 = ~n31 & n42;
  assign n44 = pi01 & ~pi05;
  assign n45 = ~n29 & n44;
  assign n46 = ~n43 & ~n45;
  assign n47 = ~n41 & ~n46;
  assign n48 = n41 & n46;
  assign n49 = ~n47 & ~n48;
  assign n50 = ~pi01 & ~n11;
  assign n51 = pi07 & ~n50;
  assign n52 = pi01 & ~n12;
  assign n53 = ~pi07 & ~n52;
  assign n54 = ~n51 & ~n53;
  assign n55 = n49 & n54;
  assign n56 = ~n49 & ~n54;
  assign n57 = ~n55 & ~n56;
  assign n58 = ~n34 & n57;
  assign n59 = n34 & ~n57;
  assign n60 = ~n58 & ~n59;
  assign n61 = ~pi01 & ~n24;
  assign n62 = pi09 & ~n61;
  assign n63 = pi01 & ~n23;
  assign n64 = ~pi09 & ~n63;
  assign n65 = ~n62 & ~n64;
  assign n66 = n60 & n65;
  assign n67 = ~n60 & ~n65;
  assign n68 = ~n66 & ~n67;
  assign n69 = n26 & n68;
  assign n70 = ~n26 & ~n68;
  assign n71 = ~n69 & ~n70;
  assign n72 = ~n58 & ~n66;
  assign n73 = ~n47 & ~n55;
  assign n74 = ~n72 & ~n73;
  assign n75 = n72 & n73;
  assign n76 = ~n74 & ~n75;
  assign n77 = n69 & ~n76;
  assign n78 = n72 & ~n73;
  assign n79 = ~n72 & n73;
  assign n80 = ~n78 & ~n79;
  assign n81 = ~n69 & ~n80;
  assign n82 = ~n77 & ~n81;
  assign po0 = n28;
  assign po1 = n71;
  assign po2 = ~n82;
endmodule
