module mul_i12_o12(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11;
  wire n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236;
  assign n13 = pi00 & pi06;
  assign n14 = pi01 & pi07;
  assign n15 = n13 & n14;
  assign n16 = pi01 & pi06;
  assign n17 = pi00 & pi07;
  assign n18 = ~n16 & ~n17;
  assign n19 = ~n15 & ~n18;
  assign n20 = pi00 & pi08;
  assign n21 = pi02 & pi06;
  assign n22 = n14 & n21;
  assign n23 = ~n14 & ~n21;
  assign n24 = ~n22 & ~n23;
  assign n25 = n20 & n24;
  assign n26 = ~n20 & ~n24;
  assign n27 = ~n25 & ~n26;
  assign n28 = n15 & n27;
  assign n29 = ~n15 & ~n27;
  assign n30 = ~n28 & ~n29;
  assign n31 = pi00 & pi09;
  assign n32 = ~n22 & ~n25;
  assign n33 = pi01 & pi08;
  assign n34 = pi03 & pi07;
  assign n35 = n21 & n34;
  assign n36 = pi03 & pi06;
  assign n37 = pi02 & pi07;
  assign n38 = ~n36 & ~n37;
  assign n39 = ~n35 & ~n38;
  assign n40 = n33 & n39;
  assign n41 = ~n33 & ~n39;
  assign n42 = ~n40 & ~n41;
  assign n43 = ~n32 & n42;
  assign n44 = n32 & ~n42;
  assign n45 = ~n43 & ~n44;
  assign n46 = n31 & n45;
  assign n47 = ~n31 & ~n45;
  assign n48 = ~n46 & ~n47;
  assign n49 = n28 & n48;
  assign n50 = ~n28 & ~n48;
  assign n51 = ~n49 & ~n50;
  assign n52 = ~n43 & ~n46;
  assign n53 = pi01 & pi10;
  assign n54 = n31 & n53;
  assign n55 = pi01 & pi09;
  assign n56 = pi00 & pi10;
  assign n57 = ~n55 & ~n56;
  assign n58 = ~n54 & ~n57;
  assign n59 = ~n35 & ~n40;
  assign n60 = pi02 & pi08;
  assign n61 = pi04 & pi06;
  assign n62 = n34 & n61;
  assign n63 = ~n34 & ~n61;
  assign n64 = ~n62 & ~n63;
  assign n65 = n60 & n64;
  assign n66 = ~n60 & ~n64;
  assign n67 = ~n65 & ~n66;
  assign n68 = ~n59 & n67;
  assign n69 = n59 & ~n67;
  assign n70 = ~n68 & ~n69;
  assign n71 = n58 & n70;
  assign n72 = ~n58 & ~n70;
  assign n73 = ~n71 & ~n72;
  assign n74 = ~n52 & n73;
  assign n75 = n52 & ~n73;
  assign n76 = ~n74 & ~n75;
  assign n77 = n49 & n76;
  assign n78 = ~n49 & ~n76;
  assign n79 = ~n77 & ~n78;
  assign n80 = ~n68 & ~n71;
  assign n81 = ~n62 & ~n65;
  assign n82 = pi03 & pi08;
  assign n83 = pi05 & pi07;
  assign n84 = n61 & n83;
  assign n85 = pi04 & pi07;
  assign n86 = pi05 & pi06;
  assign n87 = ~n85 & ~n86;
  assign n88 = ~n84 & ~n87;
  assign n89 = n82 & n88;
  assign n90 = ~n82 & ~n88;
  assign n91 = ~n89 & ~n90;
  assign n92 = ~n81 & n91;
  assign n93 = n81 & ~n91;
  assign n94 = ~n92 & ~n93;
  assign n95 = pi00 & pi11;
  assign n96 = pi02 & pi09;
  assign n97 = n53 & n96;
  assign n98 = ~n53 & ~n96;
  assign n99 = ~n97 & ~n98;
  assign n100 = n95 & n99;
  assign n101 = ~n95 & ~n99;
  assign n102 = ~n100 & ~n101;
  assign n103 = n94 & n102;
  assign n104 = ~n94 & ~n102;
  assign n105 = ~n103 & ~n104;
  assign n106 = ~n80 & n105;
  assign n107 = n80 & ~n105;
  assign n108 = ~n106 & ~n107;
  assign n109 = n54 & n108;
  assign n110 = ~n54 & ~n108;
  assign n111 = ~n109 & ~n110;
  assign n112 = n74 & n111;
  assign n113 = ~n74 & ~n111;
  assign n114 = ~n112 & ~n113;
  assign n115 = n77 & n114;
  assign n116 = ~n77 & ~n114;
  assign n117 = ~n115 & ~n116;
  assign n118 = ~n112 & ~n115;
  assign n119 = ~n106 & ~n109;
  assign n120 = ~n97 & ~n100;
  assign n121 = ~n92 & ~n103;
  assign n122 = pi05 & pi08;
  assign n123 = n85 & n122;
  assign n124 = pi04 & pi08;
  assign n125 = ~n83 & ~n124;
  assign n126 = ~n123 & ~n125;
  assign n127 = ~n84 & ~n89;
  assign n128 = n126 & ~n127;
  assign n129 = ~n126 & n127;
  assign n130 = ~n128 & ~n129;
  assign n131 = pi01 & pi11;
  assign n132 = pi03 & pi09;
  assign n133 = pi02 & pi10;
  assign n134 = ~n132 & ~n133;
  assign n135 = pi03 & pi10;
  assign n136 = n96 & n135;
  assign n137 = ~n134 & ~n136;
  assign n138 = n131 & n137;
  assign n139 = ~n131 & ~n137;
  assign n140 = ~n138 & ~n139;
  assign n141 = n130 & n140;
  assign n142 = ~n130 & ~n140;
  assign n143 = ~n141 & ~n142;
  assign n144 = ~n121 & n143;
  assign n145 = n121 & ~n143;
  assign n146 = ~n144 & ~n145;
  assign n147 = ~n120 & n146;
  assign n148 = n120 & ~n146;
  assign n149 = ~n147 & ~n148;
  assign n150 = ~n119 & n149;
  assign n151 = n119 & ~n149;
  assign n152 = ~n150 & ~n151;
  assign n153 = ~n118 & n152;
  assign n154 = n118 & ~n152;
  assign n155 = ~n153 & ~n154;
  assign n156 = ~n150 & ~n153;
  assign n157 = ~n144 & ~n147;
  assign n158 = ~n136 & ~n138;
  assign n159 = ~n128 & ~n141;
  assign n160 = ~n85 & n122;
  assign n161 = pi04 & pi09;
  assign n162 = ~n135 & ~n161;
  assign n163 = pi04 & pi10;
  assign n164 = n132 & n163;
  assign n165 = ~n162 & ~n164;
  assign n166 = pi02 & pi11;
  assign n167 = n165 & n166;
  assign n168 = ~n165 & ~n166;
  assign n169 = ~n167 & ~n168;
  assign n170 = n160 & n169;
  assign n171 = ~n160 & ~n169;
  assign n172 = ~n170 & ~n171;
  assign n173 = ~n159 & n172;
  assign n174 = n159 & ~n172;
  assign n175 = ~n173 & ~n174;
  assign n176 = ~n158 & n175;
  assign n177 = n158 & ~n175;
  assign n178 = ~n176 & ~n177;
  assign n179 = ~n157 & n178;
  assign n180 = n157 & ~n178;
  assign n181 = ~n179 & ~n180;
  assign n182 = ~n156 & n181;
  assign n183 = n156 & ~n181;
  assign n184 = ~n182 & ~n183;
  assign n185 = ~n179 & ~n182;
  assign n186 = ~n173 & ~n176;
  assign n187 = ~n164 & ~n167;
  assign n188 = ~n123 & ~n170;
  assign n189 = pi03 & pi11;
  assign n190 = pi05 & pi09;
  assign n191 = n163 & n190;
  assign n192 = ~n163 & ~n190;
  assign n193 = ~n191 & ~n192;
  assign n194 = n189 & n193;
  assign n195 = ~n189 & ~n193;
  assign n196 = ~n194 & ~n195;
  assign n197 = ~n188 & n196;
  assign n198 = n188 & ~n196;
  assign n199 = ~n197 & ~n198;
  assign n200 = ~n187 & n199;
  assign n201 = n187 & ~n199;
  assign n202 = ~n200 & ~n201;
  assign n203 = ~n186 & n202;
  assign n204 = n186 & ~n202;
  assign n205 = ~n203 & ~n204;
  assign n206 = ~n185 & n205;
  assign n207 = n185 & ~n205;
  assign n208 = ~n206 & ~n207;
  assign n209 = ~n203 & ~n206;
  assign n210 = ~n197 & ~n200;
  assign n211 = pi05 & pi11;
  assign n212 = n163 & n211;
  assign n213 = pi05 & pi10;
  assign n214 = pi04 & pi11;
  assign n215 = ~n213 & ~n214;
  assign n216 = ~n212 & ~n215;
  assign n217 = ~n191 & ~n194;
  assign n218 = n216 & ~n217;
  assign n219 = ~n216 & n217;
  assign n220 = ~n218 & ~n219;
  assign n221 = ~n210 & n220;
  assign n222 = n210 & ~n220;
  assign n223 = ~n221 & ~n222;
  assign n224 = ~n209 & n223;
  assign n225 = n209 & ~n223;
  assign n226 = ~n224 & ~n225;
  assign n227 = ~n221 & ~n224;
  assign n228 = ~n163 & n211;
  assign n229 = n218 & n228;
  assign n230 = ~n218 & ~n228;
  assign n231 = ~n229 & ~n230;
  assign n232 = ~n227 & n231;
  assign n233 = n227 & ~n231;
  assign n234 = ~n232 & ~n233;
  assign n235 = ~n212 & ~n229;
  assign n236 = ~n232 & n235;
  assign po00 = n13;
  assign po01 = n19;
  assign po02 = n30;
  assign po03 = n51;
  assign po04 = n79;
  assign po05 = n117;
  assign po06 = n155;
  assign po07 = n184;
  assign po08 = n208;
  assign po09 = n226;
  assign po10 = n234;
  assign po11 = ~n236;
endmodule
