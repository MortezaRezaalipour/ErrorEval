module mul_i12_o12 (a, b, r);
input [5:0] a, b;
output [11:0] r;


assign r = a * b;

endmodule 
