// Benchmark "circuit" written by ABC on Wed Jul 11 22:45:13 2018

module circuit ( 
    g0, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15,
    g700, g699, g698, g697, g696, g695, g694, g693, g692, g691, g690, g689,
    g688, g687, g686, g685  );
  input  g0, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14,
    g15;
  output g700, g699, g698, g697, g696, g695, g694, g693, g692, g691, g690,
    g689, g688, g687, g686, g685;
  wire g16, g17, g18, g19, g20, g21, g22, g23, g24, g25, g26, g27, g28, g29,
    g30, g31, g32, g33, g34, g35, g36, g37, g38, g39, g40, g41, g42, g43,
    g44, g45, g46, g47, g48, g49, g50, g51, g52, g53, g54, g55, g56, g57,
    g58, g59, g60, g61, g62, g63, g64, g65, g66, g67, g68, g69, g70, g71,
    g72, g73, g74, g75, g76, g77, g78, g79, g80, g81, g82, g83, g84, g85,
    g86, g87, g88, g89, g90, g91, g92, g93, g94, g95, g96, g97, g98, g99,
    g100, g101, g102, g103, g104, g105, g106, g107, g108, g109, g110, g111,
    g112, g113, g114, g115, g116, g117, g118, g119, g120, g121, g122, g123,
    g124, g125, g126, g127, g128, g129, g130, g131, g132, g133, g134, g135,
    g136, g137, g138, g139, g140, g141, g142, g143, g144, g145, g146, g147,
    g148, g149, g150, g151, g152, g153, g154, g155, g156, g157, g158, g159,
    g160, g161, g162, g163, g164, g165, g166, g167, g168, g169, g170, g171,
    g172, g173, g174, g175, g176, g177, g178, g179, g180, g181, g182, g183,
    g184, g185, g186, g187, g188, g189, g190, g191, g192, g193, g194, g195,
    g196, g197, g198, g199, g200, g201, g202, g203, g204, g205, g206, g207,
    g208, g209, g210, g211, g212, g213, g214, g215, g216, g217, g218, g219,
    g220, g221, g222, g223, g224, g225, g226, g227, g228, g229, g230, g231,
    g232, g233, g234, g235, g236, g237, g238, g239, g240, g241, g242, g243,
    g244, g245, g246, g247, g248, g249, g250, g251, g252, g253, g254, g255,
    g256, g257, g258, g259, g260, g261, g262, g263, g264, g265, g266, g267,
    g268, g269, g270, g271, g272, g273, g274, g275, g276, g277, g278, g279,
    g280, g281, g282, g283, g284, g285, g286, g287, g288, g289, g290, g291,
    g292, g293, g294, g295, g296, g297, g298, g299, g300, g301, g302, g303,
    g304, g305, g306, g307, g308, g309, g310, g311, g312, g313, g314, g315,
    g316, g317, g318, g319, g320, g321, g322, g323, g324, g325, g326, g327,
    g328, g329, g330, g331, g332, g333, g334, g335, g336, g337, g338, g339,
    g340, g341, g342, g343, g344, g345, g346, g347, g348, g349, g350, g351,
    g352, g353, g354, g355, g356, g357, g358, g359, g360, g361, g362, g363,
    g364, g365, g366, g367, g368, g369, g370, g371, g372, g373, g374, g375,
    g376, g377, g378, g379, g380, g381, g382, g383, g384, g385, g386, g387,
    g388, g389, g390, g391, g392, g393, g394, g395, g396, g397, g398, g399,
    g400, g401, g419, g420, g421, g422, g423, g424, g425, g426, g427, g428,
    g429, g430, g431, g432, g433, g434, g435, g436, g437, g438, g439, g440,
    g441, g442, g443, g444, g445, g446, g447, g448, g449, g450, g451, g452,
    g453, g454, g455, g456, g457, g458, g459, g460, g461, g462, g463, g464,
    g465, g466, g467, g468, g469, g470, g471, g472, g473, g474, g475, g476,
    g477, g478, g479, g480, g481, g482, g483, g484, g485, g486, g487, g488,
    g489, g490, g491, g492, g493, g494, g495, g496, g497, g498, g499, g500,
    g501, g502, g503, g504, g505, g506, g507, g508, g509, g510, g511, g512,
    g513, g514, g515, g516, g517, g518, g519, g520, g521, g522, g523, g524,
    g525, g526, g527, g528, g529, g530, g531, g532, g533, g534, g535, g536,
    g537, g538, g539, g540, g541, g542, g543, g544, g545, g546, g547, g548,
    g549, g550, g551, g552, g553, g554, g555, g556, g557, g558, g559, g560,
    g561, g562, g563, g564, g565, g566, g567, g568, g569, g570, g571, g572,
    g573, g574, g575, g576, g577, g578, g579, g580, g581, g582, g583, g584,
    g585, g586, g587, g588, g589, g590, g591, g592, g593, g594, g595, g596,
    g597, g598, g599, g600, g601, g602, g603, g604, g605, g606, g607, g608,
    g609, g610, g611, g612, g613, g614, g615, g616, g617, g618, g619, g620,
    g621, g622, g623, g624, g625, g626, g627, g628, g629, g630, g631, g632,
    g633, g634, g635, g636, g637, g638, g639, g648, g649, g653, g654, g655,
    g656, g657, g658, g659, g660, g661, g662, g663, g664, g665, g666, g667,
    g668, g672, g674, g675, g676, g677, g678, g679, g680, g681, g682, g683,
    g684, \0 ;
  assign g16 = g5 & g9;
  assign g17 = g7 & g8;
  assign g18 = g3 & g12;
  assign g19 = g17 & g18;
  assign g20 = g6 & g9;
  assign g21 = ~g18;
  assign g22 = g17 & g21;
  assign g23 = ~g17;
  assign g24 = g18 & g23;
  assign g25 = g22 | g24;
  assign g26 = g20 & g25;
  assign g27 = g19 | g26;
  assign g28 = g16 & g27;
  assign g29 = ~g28;
  assign g30 = g16 | g27;
  assign g31 = g29 & g30;
  assign g32 = g6 & g8;
  assign g33 = g2 & g12;
  assign g34 = ~g33;
  assign g35 = g32 & g34;
  assign g36 = ~g32;
  assign g37 = g33 & g36;
  assign g38 = g35 | g37;
  assign g39 = ~g38;
  assign g40 = g4 & g10;
  assign g41 = g39 & g40;
  assign g42 = ~g40;
  assign g43 = g38 & g42;
  assign g44 = g41 | g43;
  assign g45 = g31 & g44;
  assign g46 = g28 | g45;
  assign g47 = ~g46;
  assign g48 = g3 & g10;
  assign g49 = g32 & g33;
  assign g50 = g38 & g40;
  assign g51 = g49 | g50;
  assign g52 = g48 & g51;
  assign g53 = ~g52;
  assign g54 = g48 | g51;
  assign g55 = g53 & g54;
  assign g56 = g2 & g11;
  assign g57 = g4 & g9;
  assign g58 = ~g57;
  assign g59 = g56 & g58;
  assign g60 = ~g56;
  assign g61 = g57 & g60;
  assign g62 = g59 | g61;
  assign g63 = ~g62;
  assign g64 = g1 & g12;
  assign g65 = g63 & g64;
  assign g66 = ~g64;
  assign g67 = g62 & g66;
  assign g68 = g65 | g67;
  assign g69 = g55 & g68;
  assign g70 = ~g69;
  assign g71 = g55 | g68;
  assign g72 = g70 & g71;
  assign g73 = g5 & g8;
  assign g74 = g1 & g13;
  assign g75 = g1 & g14;
  assign g76 = g2 & g14;
  assign g77 = g3 & g14;
  assign g78 = g4 & g14;
  assign g79 = g5 & g14;
  assign g80 = g7 & g12;
  assign g81 = g79 & g80;
  assign g82 = g78 & g81;
  assign g83 = g77 & g82;
  assign g84 = g76 & g83;
  assign g85 = g75 & g84;
  assign g86 = g74 & g85;
  assign g87 = ~g86;
  assign g88 = g73 & g87;
  assign g89 = ~g73;
  assign g90 = g86 & g89;
  assign g91 = g88 | g90;
  assign g92 = ~g91;
  assign g93 = g0 & g13;
  assign g94 = g92 & g93;
  assign g95 = ~g93;
  assign g96 = g91 & g95;
  assign g97 = g94 | g96;
  assign g98 = g72 & g97;
  assign g99 = ~g98;
  assign g100 = g72 | g97;
  assign g101 = g99 & g100;
  assign g102 = g47 & g101;
  assign g103 = ~g101;
  assign g104 = g46 & g103;
  assign g105 = g102 | g104;
  assign g106 = g3 & g11;
  assign g107 = ~g85;
  assign g108 = g74 & g107;
  assign g109 = ~g74;
  assign g110 = g85 & g109;
  assign g111 = g108 | g110;
  assign g112 = g106 & g111;
  assign g113 = g0 & g14;
  assign g114 = ~g111;
  assign g115 = g106 & g114;
  assign g116 = ~g106;
  assign g117 = g111 & g116;
  assign g118 = g115 | g117;
  assign g119 = g113 & g118;
  assign g120 = g112 | g119;
  assign g121 = ~g120;
  assign g122 = ~g45;
  assign g123 = g31 | g44;
  assign g124 = g122 & g123;
  assign g125 = g5 & g10;
  assign g126 = g4 & g11;
  assign g127 = g125 & g126;
  assign g128 = ~g126;
  assign g129 = g125 & g128;
  assign g130 = ~g125;
  assign g131 = g126 & g130;
  assign g132 = g129 | g131;
  assign g133 = g7 & g9;
  assign g134 = g6 & g10;
  assign g135 = g133 & g134;
  assign g136 = g4 & g12;
  assign g137 = ~g134;
  assign g138 = g133 & g137;
  assign g139 = ~g133;
  assign g140 = g134 & g139;
  assign g141 = g138 | g140;
  assign g142 = g136 & g141;
  assign g143 = g135 | g142;
  assign g144 = g132 & g143;
  assign g145 = g127 | g144;
  assign g146 = g124 & g145;
  assign g147 = ~g118;
  assign g148 = g113 & g147;
  assign g149 = ~g113;
  assign g150 = g118 & g149;
  assign g151 = g148 | g150;
  assign g152 = ~g145;
  assign g153 = g124 & g152;
  assign g154 = ~g124;
  assign g155 = g145 & g154;
  assign g156 = g153 | g155;
  assign g157 = g151 & g156;
  assign g158 = g146 | g157;
  assign g159 = g121 & g158;
  assign g160 = ~g158;
  assign g161 = g120 & g160;
  assign g162 = g159 | g161;
  assign g163 = ~g162;
  assign g164 = g105 & g163;
  assign g165 = ~g105;
  assign g166 = g162 & g165;
  assign g167 = g164 | g166;
  assign g168 = ~g25;
  assign g169 = g20 & g168;
  assign g170 = ~g20;
  assign g171 = g25 & g170;
  assign g172 = g169 | g171;
  assign g173 = g5 & g11;
  assign g174 = g6 & g11;
  assign g175 = g7 & g10;
  assign g176 = g174 & g175;
  assign g177 = g5 & g12;
  assign g178 = ~g175;
  assign g179 = g174 & g178;
  assign g180 = ~g174;
  assign g181 = g175 & g180;
  assign g182 = g179 | g181;
  assign g183 = g177 & g182;
  assign g184 = g176 | g183;
  assign g185 = g173 & g184;
  assign g186 = ~g185;
  assign g187 = g173 | g184;
  assign g188 = g186 & g187;
  assign g189 = ~g141;
  assign g190 = g136 & g189;
  assign g191 = ~g136;
  assign g192 = g141 & g191;
  assign g193 = g190 | g192;
  assign g194 = g188 & g193;
  assign g195 = g185 | g194;
  assign g196 = g172 & g195;
  assign g197 = ~g75;
  assign g198 = g84 & g197;
  assign g199 = ~g84;
  assign g200 = g75 & g199;
  assign g201 = g198 | g200;
  assign g202 = ~g201;
  assign g203 = g2 & g13;
  assign g204 = g202 & g203;
  assign g205 = ~g203;
  assign g206 = g201 & g205;
  assign g207 = g204 | g206;
  assign g208 = ~g207;
  assign g209 = g0 & g15;
  assign g210 = g208 & g209;
  assign g211 = ~g209;
  assign g212 = g207 & g211;
  assign g213 = g210 | g212;
  assign g214 = g172 | g195;
  assign g215 = ~g196;
  assign g216 = g214 & g215;
  assign g217 = g213 & g216;
  assign g218 = g196 | g217;
  assign g219 = g201 & g203;
  assign g220 = g207 & g209;
  assign g221 = g219 | g220;
  assign g222 = g218 & g221;
  assign g223 = ~g221;
  assign g224 = g218 & g223;
  assign g225 = ~g218;
  assign g226 = g221 & g225;
  assign g227 = g224 | g226;
  assign g228 = g132 | g143;
  assign g229 = ~g144;
  assign g230 = g228 & g229;
  assign g231 = g3 & g13;
  assign g232 = ~g76;
  assign g233 = g83 & g232;
  assign g234 = ~g83;
  assign g235 = g76 & g234;
  assign g236 = g233 | g235;
  assign g237 = g231 & g236;
  assign g238 = g1 & g15;
  assign g239 = ~g236;
  assign g240 = g231 & g239;
  assign g241 = ~g231;
  assign g242 = g236 & g241;
  assign g243 = g240 | g242;
  assign g244 = g238 & g243;
  assign g245 = g237 | g244;
  assign g246 = g230 & g245;
  assign g247 = ~g245;
  assign g248 = g230 & g247;
  assign g249 = ~g230;
  assign g250 = g245 & g249;
  assign g251 = g248 | g250;
  assign g252 = ~g243;
  assign g253 = g238 & g252;
  assign g254 = ~g238;
  assign g255 = g243 & g254;
  assign g256 = g253 | g255;
  assign g257 = g4 & g13;
  assign g258 = ~g77;
  assign g259 = g82 & g258;
  assign g260 = ~g82;
  assign g261 = g77 & g260;
  assign g262 = g259 | g261;
  assign g263 = g257 & g262;
  assign g264 = g2 & g15;
  assign g265 = ~g262;
  assign g266 = g257 & g265;
  assign g267 = ~g257;
  assign g268 = g262 & g267;
  assign g269 = g266 | g268;
  assign g270 = g264 & g269;
  assign g271 = g263 | g270;
  assign g272 = g256 & g271;
  assign g273 = g256 | g271;
  assign g274 = ~g272;
  assign g275 = g273 & g274;
  assign g276 = ~g194;
  assign g277 = g188 | g193;
  assign g278 = g276 & g277;
  assign g279 = g275 & g278;
  assign g280 = g272 | g279;
  assign g281 = g251 & g280;
  assign g282 = g246 | g281;
  assign g283 = g227 & g282;
  assign g284 = g222 | g283;
  assign g285 = g167 & g284;
  assign g286 = g167 | g284;
  assign g287 = ~g285;
  assign g288 = g286 & g287;
  assign g289 = ~g151;
  assign g290 = g156 & g289;
  assign g291 = ~g156;
  assign g292 = g151 & g291;
  assign g293 = g290 | g292;
  assign g294 = g227 | g282;
  assign g295 = ~g283;
  assign g296 = g294 & g295;
  assign g297 = g293 & g296;
  assign g298 = ~g297;
  assign g299 = g293 | g296;
  assign g300 = g298 & g299;
  assign g301 = ~g217;
  assign g302 = g213 | g216;
  assign g303 = g301 & g302;
  assign g304 = g251 | g280;
  assign g305 = ~g281;
  assign g306 = g304 & g305;
  assign g307 = g303 & g306;
  assign g308 = ~g278;
  assign g309 = g275 & g308;
  assign g310 = ~g275;
  assign g311 = g278 & g310;
  assign g312 = g309 | g311;
  assign g313 = ~g182;
  assign g314 = g177 & g313;
  assign g315 = ~g177;
  assign g316 = g182 & g315;
  assign g317 = g314 | g316;
  assign g318 = g7 & g11;
  assign g319 = g6 & g12;
  assign g320 = g318 & g319;
  assign g321 = ~g319;
  assign g322 = g318 & g321;
  assign g323 = ~g318;
  assign g324 = g319 & g323;
  assign g325 = g322 | g324;
  assign g326 = g6 & g13;
  assign g327 = ~g326;
  assign g328 = g4 & g15;
  assign g329 = ~g328;
  assign g330 = g327 | g329;
  assign g331 = g7 & g13;
  assign g332 = g6 & g14;
  assign g333 = g331 & g332;
  assign g334 = ~g333;
  assign g335 = g330 & g334;
  assign g336 = ~g335;
  assign g337 = g325 & g336;
  assign g338 = g320 | g337;
  assign g339 = g317 & g338;
  assign g340 = g317 | g338;
  assign g341 = ~g339;
  assign g342 = g340 & g341;
  assign g343 = g5 & g13;
  assign g344 = ~g78;
  assign g345 = g81 & g344;
  assign g346 = ~g81;
  assign g347 = g78 & g346;
  assign g348 = g345 | g347;
  assign g349 = g343 & g348;
  assign g350 = g3 & g15;
  assign g351 = ~g348;
  assign g352 = g343 & g351;
  assign g353 = ~g343;
  assign g354 = g348 & g353;
  assign g355 = g352 | g354;
  assign g356 = g350 & g355;
  assign g357 = g349 | g356;
  assign g358 = g342 & g357;
  assign g359 = g339 | g358;
  assign g360 = g312 & g359;
  assign g361 = g312 | g359;
  assign g362 = ~g360;
  assign g363 = g361 & g362;
  assign g364 = ~g357;
  assign g365 = g342 & g364;
  assign g366 = ~g342;
  assign g367 = g357 & g366;
  assign g368 = g365 | g367;
  assign g369 = ~g269;
  assign g370 = g264 & g369;
  assign g371 = ~g264;
  assign g372 = g269 & g371;
  assign g373 = g370 | g372;
  assign g374 = g368 & g373;
  assign g375 = ~g355;
  assign g376 = g350 & g375;
  assign g377 = ~g350;
  assign g378 = g355 & g377;
  assign g379 = g376 | g378;
  assign g380 = ~g325;
  assign g381 = g335 & g380;
  assign g382 = g337 | g381;
  assign g383 = ~g382;
  assign g384 = g379 & g383;
  assign g385 = ~g379;
  assign g386 = g382 & g385;
  assign g387 = g384 | g386;
  assign g388 = ~g387;
  assign g389 = g326 & g329;
  assign g390 = g327 & g328;
  assign g391 = g389 | g390;
  assign g392 = ~g391;
  assign g393 = g333 & g392;
  assign g394 = g334 & g391;
  assign g395 = g393 | g394;
  assign g396 = ~g79;
  assign g397 = g80 & g396;
  assign g398 = ~g80;
  assign g399 = g79 & g398;
  assign g400 = g397 | g399;
  assign g401 = g395 & g400;
  assign g419 = ~g395;
  assign g420 = g400 & g419;
  assign g421 = ~g400;
  assign g422 = g395 & g421;
  assign g423 = g420 | g422;
  assign g424 = \0  & g423;
  assign g425 = g401 | g424;
  assign g426 = g388 & g425;
  assign g427 = g384 | g426;
  assign g428 = ~g368;
  assign g429 = g373 & g428;
  assign g430 = ~g373;
  assign g431 = g368 & g430;
  assign g432 = g429 | g431;
  assign g433 = g427 & g432;
  assign g434 = g374 | g433;
  assign g435 = g363 & g434;
  assign g436 = g360 | g435;
  assign g437 = ~g306;
  assign g438 = g303 & g437;
  assign g439 = ~g303;
  assign g440 = g306 & g439;
  assign g441 = g438 | g440;
  assign g442 = g436 & g441;
  assign g443 = g307 | g442;
  assign g444 = g300 & g443;
  assign g445 = g297 | g444;
  assign g446 = g288 & g445;
  assign g447 = g285 | g446;
  assign g448 = ~g447;
  assign g449 = g120 & g158;
  assign g450 = g105 & g162;
  assign g451 = g449 | g450;
  assign g452 = g52 | g69;
  assign g453 = g4 & g8;
  assign g454 = g0 & g12;
  assign g455 = ~g454;
  assign g456 = g453 & g455;
  assign g457 = ~g453;
  assign g458 = g454 & g457;
  assign g459 = g456 | g458;
  assign g460 = ~g459;
  assign g461 = g3 & g9;
  assign g462 = g460 & g461;
  assign g463 = ~g461;
  assign g464 = g459 & g463;
  assign g465 = g462 | g464;
  assign g466 = g452 | g465;
  assign g467 = g452 & g465;
  assign g468 = ~g467;
  assign g469 = g466 & g468;
  assign g470 = ~g469;
  assign g471 = g56 & g57;
  assign g472 = g62 & g64;
  assign g473 = g471 | g472;
  assign g474 = g2 & g10;
  assign g475 = g1 & g11;
  assign g476 = ~g475;
  assign g477 = g474 & g476;
  assign g478 = ~g474;
  assign g479 = g475 & g478;
  assign g480 = g477 | g479;
  assign g481 = g473 | g480;
  assign g482 = g473 & g480;
  assign g483 = ~g482;
  assign g484 = g481 & g483;
  assign g485 = g470 & g484;
  assign g486 = ~g484;
  assign g487 = g469 & g486;
  assign g488 = g485 | g487;
  assign g489 = g73 & g86;
  assign g490 = g91 & g93;
  assign g491 = g489 | g490;
  assign g492 = ~g491;
  assign g493 = g46 & g101;
  assign g494 = g98 | g493;
  assign g495 = g492 & g494;
  assign g496 = ~g494;
  assign g497 = g491 & g496;
  assign g498 = g495 | g497;
  assign g499 = ~g498;
  assign g500 = g488 & g499;
  assign g501 = ~g488;
  assign g502 = g498 & g501;
  assign g503 = g500 | g502;
  assign g504 = g451 | g503;
  assign g505 = g451 & g503;
  assign g506 = ~g505;
  assign g507 = g504 & g506;
  assign g508 = g448 & g507;
  assign g509 = ~g507;
  assign g510 = g447 & g509;
  assign g511 = g447 & g507;
  assign g512 = g505 | g511;
  assign g513 = g491 & g494;
  assign g514 = g488 & g498;
  assign g515 = g513 | g514;
  assign g516 = ~g515;
  assign g517 = g469 & g484;
  assign g518 = g467 | g517;
  assign g519 = g474 & g475;
  assign g520 = g482 | g519;
  assign g521 = ~g520;
  assign g522 = g3 & g8;
  assign g523 = g0 & g11;
  assign g524 = ~g523;
  assign g525 = g522 & g524;
  assign g526 = ~g522;
  assign g527 = g523 & g526;
  assign g528 = g525 | g527;
  assign g529 = ~g528;
  assign g530 = g1 & g10;
  assign g531 = g529 & g530;
  assign g532 = ~g530;
  assign g533 = g528 & g532;
  assign g534 = g531 | g533;
  assign g535 = g2 & g9;
  assign g536 = g453 & g454;
  assign g537 = g459 & g461;
  assign g538 = g536 | g537;
  assign g539 = g535 & g538;
  assign g540 = ~g539;
  assign g541 = g535 | g538;
  assign g542 = g540 & g541;
  assign g543 = g534 & g542;
  assign g544 = ~g543;
  assign g545 = g534 | g542;
  assign g546 = g544 & g545;
  assign g547 = g521 & g546;
  assign g548 = ~g546;
  assign g549 = g520 & g548;
  assign g550 = g547 | g549;
  assign g551 = g518 | g550;
  assign g552 = g518 & g550;
  assign g553 = ~g552;
  assign g554 = g551 & g553;
  assign g555 = g516 & g554;
  assign g556 = ~g554;
  assign g557 = g515 & g556;
  assign g558 = g555 | g557;
  assign g559 = g512 & g558;
  assign g560 = ~g559;
  assign g561 = g512 | g558;
  assign g562 = g515 & g554;
  assign g563 = g559 | g562;
  assign g564 = ~g563;
  assign g565 = g520 & g546;
  assign g566 = g552 | g565;
  assign g567 = g539 | g543;
  assign g568 = ~g567;
  assign g569 = g522 & g523;
  assign g570 = g528 & g530;
  assign g571 = g569 | g570;
  assign g572 = g2 & g8;
  assign g573 = g0 & g10;
  assign g574 = ~g573;
  assign g575 = g572 & g574;
  assign g576 = ~g572;
  assign g577 = g573 & g576;
  assign g578 = g575 | g577;
  assign g579 = ~g578;
  assign g580 = g1 & g9;
  assign g581 = g579 & g580;
  assign g582 = ~g580;
  assign g583 = g578 & g582;
  assign g584 = g581 | g583;
  assign g585 = g571 | g584;
  assign g586 = g571 & g584;
  assign g587 = ~g586;
  assign g588 = g585 & g587;
  assign g589 = g568 & g588;
  assign g590 = ~g588;
  assign g591 = g567 & g590;
  assign g592 = g589 | g591;
  assign g593 = g566 | g592;
  assign g594 = g566 & g592;
  assign g595 = ~g594;
  assign g596 = g593 & g595;
  assign g597 = g564 & g596;
  assign g598 = ~g596;
  assign g599 = g563 & g598;
  assign g600 = g563 & g596;
  assign g601 = g594 | g600;
  assign g602 = g567 & g588;
  assign g603 = g586 | g602;
  assign g604 = ~g603;
  assign g605 = g572 & g573;
  assign g606 = g578 & g580;
  assign g607 = g605 | g606;
  assign g608 = g1 & g8;
  assign g609 = g0 & g9;
  assign g610 = ~g609;
  assign g611 = g608 & g610;
  assign g612 = ~g608;
  assign g613 = g609 & g612;
  assign g614 = g611 | g613;
  assign g615 = g607 | g614;
  assign g616 = g607 & g614;
  assign g617 = ~g616;
  assign g618 = g615 & g617;
  assign g619 = g604 & g618;
  assign g620 = ~g618;
  assign g621 = g603 & g620;
  assign g622 = g619 | g621;
  assign g623 = g601 & g622;
  assign g624 = ~g623;
  assign g625 = g601 | g622;
  assign g626 = g603 & g618;
  assign g627 = g623 | g626;
  assign g628 = ~g627;
  assign g629 = g0 & g8;
  assign g630 = g608 & g609;
  assign g631 = g616 | g630;
  assign g632 = g629 & g631;
  assign g633 = ~g632;
  assign g634 = g629 | g631;
  assign g635 = g633 & g634;
  assign g636 = g628 & g635;
  assign g637 = ~g635;
  assign g638 = g627 & g637;
  assign g639 = g627 & g635;
  assign g648 = ~g424;
  assign g649 = \0  | g423;
  assign g653 = ~g433;
  assign g654 = g427 | g432;
  assign g655 = ~g434;
  assign g656 = g363 & g655;
  assign g657 = ~g363;
  assign g658 = g434 & g657;
  assign g659 = ~g442;
  assign g660 = g436 | g441;
  assign g661 = ~g443;
  assign g662 = g300 & g661;
  assign g663 = ~g300;
  assign g664 = g443 & g663;
  assign g665 = ~g445;
  assign g666 = g288 & g665;
  assign g667 = ~g288;
  assign g668 = g445 & g667;
  assign g672 = g648 & g649;
  assign g674 = g653 & g654;
  assign g675 = g656 | g658;
  assign g676 = g659 & g660;
  assign g677 = g662 | g664;
  assign g678 = g666 | g668;
  assign g679 = g508 | g510;
  assign g680 = g560 & g561;
  assign g681 = g597 | g599;
  assign g682 = g624 & g625;
  assign g683 = g636 | g638;
  assign g684 = g632 | g639;
  assign g685 = \0 ;
  assign g686 = \0 ;
  assign g687 = \0 ;
  assign g688 = g672;
  assign g689 = \0 ;
  assign g690 = g674;
  assign g691 = g675;
  assign g692 = g676;
  assign g693 = g677;
  assign g694 = g678;
  assign g695 = g679;
  assign g696 = g680;
  assign g697 = g681;
  assign g698 = g682;
  assign g699 = g683;
  assign g700 = g684;
  assign \0  = 1'b0;
endmodule


