module adder_i8_o5(pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, po0, po1, po2, po3, po4);
  input pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7;
  output po0, po1, po2, po3, po4;
  wire n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32;
  assign n9 = pi0 & pi4;
  assign n10 = ~pi0 & ~pi4;
  assign n11 = ~n9 & ~n10;
  assign n12 = pi1 & pi5;
  assign n13 = ~pi1 & ~pi5;
  assign n14 = ~n12 & ~n13;
  assign n15 = n9 & n14;
  assign n16 = ~n9 & ~n14;
  assign n17 = ~n15 & ~n16;
  assign n18 = ~n12 & ~n15;
  assign n19 = pi2 & pi6;
  assign n20 = ~pi2 & ~pi6;
  assign n21 = ~n19 & ~n20;
  assign n22 = ~n18 & n21;
  assign n23 = n18 & ~n21;
  assign n24 = ~n22 & ~n23;
  assign n25 = ~n19 & ~n22;
  assign n26 = pi3 & pi7;
  assign n27 = ~pi3 & ~pi7;
  assign n28 = ~n26 & ~n27;
  assign n29 = ~n25 & n28;
  assign n30 = n25 & ~n28;
  assign n31 = ~n29 & ~n30;
  assign n32 = ~n26 & ~n29;
  assign po0 = n11;
  assign po1 = n17;
  assign po2 = n24;
  assign po3 = n31;
  assign po4 = ~n32;
endmodule
