module adder_i44_o23 (a,b,r);
input [21:0] a,b;
output [22:0] r;

assign r = a+b;

endmodule

