module top(pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, po0, po1, po2, po3, po4, po5, po6, po7);
  input pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93;
  assign n9 = pi0 & pi4;
  assign n10 = pi0 & pi5;
  assign n11 = pi1 & pi4;
  assign n12 = ~n10 & ~n11;
  assign n13 = n10 & n11;
  assign n14 = ~n12 & ~n13;
  assign n15 = pi2 & pi5;
  assign n16 = n11 & n15;
  assign n17 = pi1 & pi5;
  assign n18 = pi2 & pi4;
  assign n19 = ~n17 & ~n18;
  assign n20 = ~n16 & ~n19;
  assign n21 = pi0 & pi6;
  assign n22 = ~n20 & ~n21;
  assign n23 = n20 & n21;
  assign n24 = ~n22 & ~n23;
  assign n25 = n13 & n24;
  assign n26 = ~n13 & ~n24;
  assign n27 = ~n25 & ~n26;
  assign n28 = pi0 & pi7;
  assign n29 = ~n16 & ~n23;
  assign n30 = pi1 & pi6;
  assign n31 = pi3 & pi4;
  assign n32 = n15 & n31;
  assign n33 = ~n15 & ~n31;
  assign n34 = ~n32 & ~n33;
  assign n35 = n30 & n34;
  assign n36 = ~n30 & ~n34;
  assign n37 = ~n35 & ~n36;
  assign n38 = ~n29 & n37;
  assign n39 = n29 & ~n37;
  assign n40 = ~n38 & ~n39;
  assign n41 = n28 & n40;
  assign n42 = ~n28 & ~n40;
  assign n43 = ~n41 & ~n42;
  assign n44 = n25 & n43;
  assign n45 = ~n25 & ~n43;
  assign n46 = ~n44 & ~n45;
  assign n47 = ~n38 & ~n41;
  assign n48 = pi1 & pi7;
  assign n49 = pi3 & pi5;
  assign n50 = pi2 & pi6;
  assign n51 = ~n49 & ~n50;
  assign n52 = pi3 & pi6;
  assign n53 = n15 & n52;
  assign n54 = ~n51 & ~n53;
  assign n55 = ~n32 & ~n35;
  assign n56 = n54 & ~n55;
  assign n57 = ~n54 & n55;
  assign n58 = ~n56 & ~n57;
  assign n59 = n48 & n58;
  assign n60 = ~n48 & ~n58;
  assign n61 = ~n59 & ~n60;
  assign n62 = ~n47 & n61;
  assign n63 = n47 & ~n61;
  assign n64 = ~n62 & ~n63;
  assign n65 = n44 & n64;
  assign n66 = ~n44 & ~n64;
  assign n67 = ~n65 & ~n66;
  assign n68 = ~n62 & ~n65;
  assign n69 = ~n56 & ~n59;
  assign n70 = pi2 & pi7;
  assign n71 = ~n15 & n52;
  assign n72 = n70 & n71;
  assign n73 = ~n70 & ~n71;
  assign n74 = ~n72 & ~n73;
  assign n75 = ~n69 & n74;
  assign n76 = n69 & ~n74;
  assign n77 = ~n75 & ~n76;
  assign n78 = n68 & n77;
  assign n79 = ~n68 & ~n77;
  assign n80 = ~n78 & ~n79;
  assign n81 = ~n53 & ~n72;
  assign n82 = pi3 & pi7;
  assign n83 = ~n81 & n82;
  assign n84 = n81 & ~n82;
  assign n85 = ~n83 & ~n84;
  assign n86 = n62 & ~n76;
  assign n87 = ~n75 & ~n86;
  assign n88 = n85 & ~n87;
  assign n89 = ~n62 & ~n75;
  assign n90 = ~n76 & ~n89;
  assign n91 = ~n85 & ~n90;
  assign n92 = ~n88 & ~n91;
  assign n93 = ~n83 & ~n88;
  assign po0 = n9;
  assign po1 = n14;
  assign po2 = n27;
  assign po3 = n46;
  assign po4 = n67;
  assign po5 = ~n80;
  assign po6 = n92;
  assign po7 = ~n93;
endmodule
