module adder_i20_o11 (a,b,r);
input [9:0] a,b;
output [10:0] r;

assign r = a+b;

endmodule

