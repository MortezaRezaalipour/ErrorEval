module adder_i32_o17 (a,b,r);
input [15:0] a,b;
output [16:0] r;

assign r = a+b;

endmodule

