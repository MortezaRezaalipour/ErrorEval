module top(pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, po0, po1, po2, po3);
  input pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7;
  output po0, po1, po2, po3;
  wire n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52;
  assign n9 = pi0 & ~pi4;
  assign n10 = ~pi0 & pi4;
  assign n11 = ~n9 & ~n10;
  assign n12 = ~pi1 & pi5;
  assign n13 = pi1 & ~pi5;
  assign n14 = ~n12 & ~n13;
  assign n15 = pi3 & ~pi7;
  assign n16 = ~pi3 & pi7;
  assign n17 = ~pi2 & pi6;
  assign n18 = pi2 & ~pi6;
  assign n19 = ~n9 & ~n13;
  assign n20 = ~n12 & ~n19;
  assign n21 = ~n18 & ~n20;
  assign n22 = ~n17 & ~n21;
  assign n23 = ~n16 & n22;
  assign n24 = ~n15 & ~n23;
  assign n25 = ~n10 & ~n24;
  assign n26 = ~n15 & ~n22;
  assign n27 = ~n16 & ~n26;
  assign n28 = ~n9 & ~n27;
  assign n29 = ~n25 & ~n28;
  assign n30 = ~n14 & ~n29;
  assign n31 = n9 & ~n27;
  assign n32 = n10 & ~n24;
  assign n33 = ~n31 & ~n32;
  assign n34 = n14 & ~n33;
  assign n35 = ~n30 & ~n34;
  assign n36 = ~n17 & ~n18;
  assign n37 = n10 & ~n13;
  assign n38 = ~n12 & ~n37;
  assign n39 = ~n24 & n38;
  assign n40 = ~n20 & ~n27;
  assign n41 = ~n39 & ~n40;
  assign n42 = ~n36 & ~n41;
  assign n43 = n20 & ~n27;
  assign n44 = ~n24 & ~n38;
  assign n45 = ~n43 & ~n44;
  assign n46 = n36 & ~n45;
  assign n47 = ~n42 & ~n46;
  assign n48 = n16 & ~n22;
  assign n49 = ~n18 & ~n38;
  assign n50 = n15 & ~n17;
  assign n51 = ~n49 & n50;
  assign n52 = ~n48 & ~n51;
  assign po0 = ~n11;
  assign po1 = ~n35;
  assign po2 = ~n47;
  assign po3 = ~n52;
endmodule
