module top(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, po0, po1, po2, po3, po4, po5);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11;
  output po0, po1, po2, po3, po4, po5;
  wire n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89;
  assign n13 = pi00 & ~pi06;
  assign n14 = ~pi00 & pi06;
  assign n15 = ~n13 & ~n14;
  assign n16 = ~pi01 & pi07;
  assign n17 = pi01 & ~pi07;
  assign n18 = ~n16 & ~n17;
  assign n19 = pi05 & ~pi11;
  assign n20 = ~pi05 & pi11;
  assign n21 = ~pi04 & pi10;
  assign n22 = pi04 & ~pi10;
  assign n23 = ~pi03 & pi09;
  assign n24 = pi03 & ~pi09;
  assign n25 = pi02 & ~pi08;
  assign n26 = ~n24 & ~n25;
  assign n27 = ~pi02 & pi08;
  assign n28 = n13 & ~n16;
  assign n29 = ~n17 & ~n28;
  assign n30 = ~n27 & ~n29;
  assign n31 = n26 & ~n30;
  assign n32 = ~n23 & ~n31;
  assign n33 = ~n22 & ~n32;
  assign n34 = ~n21 & ~n33;
  assign n35 = ~n20 & n34;
  assign n36 = ~n19 & ~n35;
  assign n37 = ~n14 & ~n36;
  assign n38 = ~n19 & ~n34;
  assign n39 = ~n20 & ~n38;
  assign n40 = ~n13 & ~n39;
  assign n41 = ~n37 & ~n40;
  assign n42 = ~n18 & ~n41;
  assign n43 = n13 & ~n39;
  assign n44 = n14 & ~n36;
  assign n45 = ~n43 & ~n44;
  assign n46 = n18 & ~n45;
  assign n47 = ~n42 & ~n46;
  assign n48 = ~n25 & ~n27;
  assign n49 = ~n14 & ~n16;
  assign n50 = ~n17 & ~n49;
  assign n51 = ~n36 & n50;
  assign n52 = ~n29 & ~n39;
  assign n53 = ~n51 & ~n52;
  assign n54 = n48 & ~n53;
  assign n55 = n29 & ~n39;
  assign n56 = ~n36 & ~n50;
  assign n57 = ~n55 & ~n56;
  assign n58 = ~n48 & ~n57;
  assign n59 = ~n54 & ~n58;
  assign n60 = ~n23 & ~n24;
  assign n61 = ~n27 & ~n50;
  assign n62 = ~n25 & ~n61;
  assign n63 = ~n36 & ~n62;
  assign n64 = ~n25 & ~n30;
  assign n65 = ~n39 & n64;
  assign n66 = ~n63 & ~n65;
  assign n67 = ~n60 & ~n66;
  assign n68 = ~n36 & n62;
  assign n69 = ~n39 & ~n64;
  assign n70 = ~n68 & ~n69;
  assign n71 = n60 & ~n70;
  assign n72 = ~n67 & ~n71;
  assign n73 = ~n21 & ~n22;
  assign n74 = n32 & ~n39;
  assign n75 = n26 & ~n61;
  assign n76 = ~n23 & ~n75;
  assign n77 = ~n36 & ~n76;
  assign n78 = ~n74 & ~n77;
  assign n79 = n73 & ~n78;
  assign n80 = ~n36 & n76;
  assign n81 = ~n32 & ~n39;
  assign n82 = ~n80 & ~n81;
  assign n83 = ~n73 & ~n82;
  assign n84 = ~n79 & ~n83;
  assign n85 = n20 & ~n34;
  assign n86 = ~n22 & ~n76;
  assign n87 = n19 & ~n21;
  assign n88 = ~n86 & n87;
  assign n89 = ~n85 & ~n88;
  assign po0 = ~n15;
  assign po1 = ~n47;
  assign po2 = ~n59;
  assign po3 = ~n72;
  assign po4 = ~n84;
  assign po5 = ~n89;
endmodule
