module adder_i36_o19 (a,b,r);
input [17:0] a,b;
output [18:0] r;

assign r = a+b;

endmodule

