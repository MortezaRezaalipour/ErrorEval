module adder_i40_o21 (a,b,r);
input [19:0] a,b;
output [20:0] r;

assign r = a+b;

endmodule

