module sad_i10_o3(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, po0, po1, po2);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09;
  output po0, po1, po2;
  wire n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79;
  assign n11 = ~pi02 & ~pi04;
  assign n12 = pi02 & pi04;
  assign n13 = ~n11 & ~n12;
  assign n14 = ~pi00 & pi06;
  assign n15 = pi00 & ~pi06;
  assign n16 = ~n14 & ~n15;
  assign n17 = n13 & n16;
  assign n18 = ~n13 & ~n16;
  assign n19 = ~n17 & ~n18;
  assign n20 = ~pi00 & pi08;
  assign n21 = pi00 & ~pi08;
  assign n22 = ~n20 & ~n21;
  assign n23 = ~n19 & ~n22;
  assign n24 = n19 & n22;
  assign n25 = ~n23 & ~n24;
  assign n26 = pi00 & ~pi04;
  assign n27 = ~pi01 & pi05;
  assign n28 = ~n26 & n27;
  assign n29 = ~pi00 & pi04;
  assign n30 = pi01 & ~pi05;
  assign n31 = ~n29 & n30;
  assign n32 = ~n28 & ~n31;
  assign n33 = pi00 & ~pi02;
  assign n34 = ~pi01 & pi03;
  assign n35 = ~n33 & n34;
  assign n36 = ~pi00 & pi02;
  assign n37 = pi01 & ~pi03;
  assign n38 = ~n36 & n37;
  assign n39 = ~n35 & ~n38;
  assign n40 = ~n32 & ~n39;
  assign n41 = n32 & n39;
  assign n42 = ~n40 & ~n41;
  assign n43 = ~pi01 & ~n15;
  assign n44 = pi07 & ~n43;
  assign n45 = pi01 & ~n14;
  assign n46 = ~pi07 & ~n45;
  assign n47 = ~n44 & ~n46;
  assign n48 = n42 & n47;
  assign n49 = ~n42 & ~n47;
  assign n50 = ~n48 & ~n49;
  assign n51 = pi00 & ~n12;
  assign n52 = ~pi00 & ~n11;
  assign n53 = ~n51 & ~n52;
  assign n54 = ~n17 & ~n53;
  assign n55 = n50 & n54;
  assign n56 = ~n50 & ~n54;
  assign n57 = ~n55 & ~n56;
  assign n58 = ~pi01 & ~n21;
  assign n59 = pi09 & ~n58;
  assign n60 = pi01 & ~n20;
  assign n61 = ~pi09 & ~n60;
  assign n62 = ~n59 & ~n61;
  assign n63 = n57 & n62;
  assign n64 = ~n57 & ~n62;
  assign n65 = ~n63 & ~n64;
  assign n66 = n23 & n65;
  assign n67 = ~n23 & ~n65;
  assign n68 = ~n66 & ~n67;
  assign n69 = ~n40 & ~n48;
  assign n70 = ~n55 & ~n63;
  assign n71 = n69 & ~n70;
  assign n72 = ~n69 & n70;
  assign n73 = ~n71 & ~n72;
  assign n74 = ~n66 & ~n73;
  assign n75 = n69 & n70;
  assign n76 = ~n69 & ~n70;
  assign n77 = ~n75 & ~n76;
  assign n78 = n66 & ~n77;
  assign n79 = ~n74 & ~n78;
  assign po0 = n25;
  assign po1 = n68;
  assign po2 = ~n79;
endmodule
