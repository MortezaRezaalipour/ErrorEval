module adder_i8_o5_tb;
reg [7:0] pi;
wire [4:0] po;
adder_i8_o5 dut( pi[0] , pi[1] , pi[2] , pi[3] , pi[4] , pi[5] , pi[6] , pi[7] , po[0] , po[1] , po[2] , po[3] , po[4] );
initial
begin
# 1  pi=8'b00000000;
#1 $display("%b", po);
# 1  pi=8'b00000001;
#1 $display("%b", po);
# 1  pi=8'b00000010;
#1 $display("%b", po);
# 1  pi=8'b00000011;
#1 $display("%b", po);
# 1  pi=8'b00000100;
#1 $display("%b", po);
# 1  pi=8'b00000101;
#1 $display("%b", po);
# 1  pi=8'b00000110;
#1 $display("%b", po);
# 1  pi=8'b00000111;
#1 $display("%b", po);
# 1  pi=8'b00001000;
#1 $display("%b", po);
# 1  pi=8'b00001001;
#1 $display("%b", po);
# 1  pi=8'b00001010;
#1 $display("%b", po);
# 1  pi=8'b00001011;
#1 $display("%b", po);
# 1  pi=8'b00001100;
#1 $display("%b", po);
# 1  pi=8'b00001101;
#1 $display("%b", po);
# 1  pi=8'b00001110;
#1 $display("%b", po);
# 1  pi=8'b00001111;
#1 $display("%b", po);
# 1  pi=8'b00010000;
#1 $display("%b", po);
# 1  pi=8'b00010001;
#1 $display("%b", po);
# 1  pi=8'b00010010;
#1 $display("%b", po);
# 1  pi=8'b00010011;
#1 $display("%b", po);
# 1  pi=8'b00010100;
#1 $display("%b", po);
# 1  pi=8'b00010101;
#1 $display("%b", po);
# 1  pi=8'b00010110;
#1 $display("%b", po);
# 1  pi=8'b00010111;
#1 $display("%b", po);
# 1  pi=8'b00011000;
#1 $display("%b", po);
# 1  pi=8'b00011001;
#1 $display("%b", po);
# 1  pi=8'b00011010;
#1 $display("%b", po);
# 1  pi=8'b00011011;
#1 $display("%b", po);
# 1  pi=8'b00011100;
#1 $display("%b", po);
# 1  pi=8'b00011101;
#1 $display("%b", po);
# 1  pi=8'b00011110;
#1 $display("%b", po);
# 1  pi=8'b00011111;
#1 $display("%b", po);
# 1  pi=8'b00100000;
#1 $display("%b", po);
# 1  pi=8'b00100001;
#1 $display("%b", po);
# 1  pi=8'b00100010;
#1 $display("%b", po);
# 1  pi=8'b00100011;
#1 $display("%b", po);
# 1  pi=8'b00100100;
#1 $display("%b", po);
# 1  pi=8'b00100101;
#1 $display("%b", po);
# 1  pi=8'b00100110;
#1 $display("%b", po);
# 1  pi=8'b00100111;
#1 $display("%b", po);
# 1  pi=8'b00101000;
#1 $display("%b", po);
# 1  pi=8'b00101001;
#1 $display("%b", po);
# 1  pi=8'b00101010;
#1 $display("%b", po);
# 1  pi=8'b00101011;
#1 $display("%b", po);
# 1  pi=8'b00101100;
#1 $display("%b", po);
# 1  pi=8'b00101101;
#1 $display("%b", po);
# 1  pi=8'b00101110;
#1 $display("%b", po);
# 1  pi=8'b00101111;
#1 $display("%b", po);
# 1  pi=8'b00110000;
#1 $display("%b", po);
# 1  pi=8'b00110001;
#1 $display("%b", po);
# 1  pi=8'b00110010;
#1 $display("%b", po);
# 1  pi=8'b00110011;
#1 $display("%b", po);
# 1  pi=8'b00110100;
#1 $display("%b", po);
# 1  pi=8'b00110101;
#1 $display("%b", po);
# 1  pi=8'b00110110;
#1 $display("%b", po);
# 1  pi=8'b00110111;
#1 $display("%b", po);
# 1  pi=8'b00111000;
#1 $display("%b", po);
# 1  pi=8'b00111001;
#1 $display("%b", po);
# 1  pi=8'b00111010;
#1 $display("%b", po);
# 1  pi=8'b00111011;
#1 $display("%b", po);
# 1  pi=8'b00111100;
#1 $display("%b", po);
# 1  pi=8'b00111101;
#1 $display("%b", po);
# 1  pi=8'b00111110;
#1 $display("%b", po);
# 1  pi=8'b00111111;
#1 $display("%b", po);
# 1  pi=8'b01000000;
#1 $display("%b", po);
# 1  pi=8'b01000001;
#1 $display("%b", po);
# 1  pi=8'b01000010;
#1 $display("%b", po);
# 1  pi=8'b01000011;
#1 $display("%b", po);
# 1  pi=8'b01000100;
#1 $display("%b", po);
# 1  pi=8'b01000101;
#1 $display("%b", po);
# 1  pi=8'b01000110;
#1 $display("%b", po);
# 1  pi=8'b01000111;
#1 $display("%b", po);
# 1  pi=8'b01001000;
#1 $display("%b", po);
# 1  pi=8'b01001001;
#1 $display("%b", po);
# 1  pi=8'b01001010;
#1 $display("%b", po);
# 1  pi=8'b01001011;
#1 $display("%b", po);
# 1  pi=8'b01001100;
#1 $display("%b", po);
# 1  pi=8'b01001101;
#1 $display("%b", po);
# 1  pi=8'b01001110;
#1 $display("%b", po);
# 1  pi=8'b01001111;
#1 $display("%b", po);
# 1  pi=8'b01010000;
#1 $display("%b", po);
# 1  pi=8'b01010001;
#1 $display("%b", po);
# 1  pi=8'b01010010;
#1 $display("%b", po);
# 1  pi=8'b01010011;
#1 $display("%b", po);
# 1  pi=8'b01010100;
#1 $display("%b", po);
# 1  pi=8'b01010101;
#1 $display("%b", po);
# 1  pi=8'b01010110;
#1 $display("%b", po);
# 1  pi=8'b01010111;
#1 $display("%b", po);
# 1  pi=8'b01011000;
#1 $display("%b", po);
# 1  pi=8'b01011001;
#1 $display("%b", po);
# 1  pi=8'b01011010;
#1 $display("%b", po);
# 1  pi=8'b01011011;
#1 $display("%b", po);
# 1  pi=8'b01011100;
#1 $display("%b", po);
# 1  pi=8'b01011101;
#1 $display("%b", po);
# 1  pi=8'b01011110;
#1 $display("%b", po);
# 1  pi=8'b01011111;
#1 $display("%b", po);
# 1  pi=8'b01100000;
#1 $display("%b", po);
# 1  pi=8'b01100001;
#1 $display("%b", po);
# 1  pi=8'b01100010;
#1 $display("%b", po);
# 1  pi=8'b01100011;
#1 $display("%b", po);
# 1  pi=8'b01100100;
#1 $display("%b", po);
# 1  pi=8'b01100101;
#1 $display("%b", po);
# 1  pi=8'b01100110;
#1 $display("%b", po);
# 1  pi=8'b01100111;
#1 $display("%b", po);
# 1  pi=8'b01101000;
#1 $display("%b", po);
# 1  pi=8'b01101001;
#1 $display("%b", po);
# 1  pi=8'b01101010;
#1 $display("%b", po);
# 1  pi=8'b01101011;
#1 $display("%b", po);
# 1  pi=8'b01101100;
#1 $display("%b", po);
# 1  pi=8'b01101101;
#1 $display("%b", po);
# 1  pi=8'b01101110;
#1 $display("%b", po);
# 1  pi=8'b01101111;
#1 $display("%b", po);
# 1  pi=8'b01110000;
#1 $display("%b", po);
# 1  pi=8'b01110001;
#1 $display("%b", po);
# 1  pi=8'b01110010;
#1 $display("%b", po);
# 1  pi=8'b01110011;
#1 $display("%b", po);
# 1  pi=8'b01110100;
#1 $display("%b", po);
# 1  pi=8'b01110101;
#1 $display("%b", po);
# 1  pi=8'b01110110;
#1 $display("%b", po);
# 1  pi=8'b01110111;
#1 $display("%b", po);
# 1  pi=8'b01111000;
#1 $display("%b", po);
# 1  pi=8'b01111001;
#1 $display("%b", po);
# 1  pi=8'b01111010;
#1 $display("%b", po);
# 1  pi=8'b01111011;
#1 $display("%b", po);
# 1  pi=8'b01111100;
#1 $display("%b", po);
# 1  pi=8'b01111101;
#1 $display("%b", po);
# 1  pi=8'b01111110;
#1 $display("%b", po);
# 1  pi=8'b01111111;
#1 $display("%b", po);
# 1  pi=8'b10000000;
#1 $display("%b", po);
# 1  pi=8'b10000001;
#1 $display("%b", po);
# 1  pi=8'b10000010;
#1 $display("%b", po);
# 1  pi=8'b10000011;
#1 $display("%b", po);
# 1  pi=8'b10000100;
#1 $display("%b", po);
# 1  pi=8'b10000101;
#1 $display("%b", po);
# 1  pi=8'b10000110;
#1 $display("%b", po);
# 1  pi=8'b10000111;
#1 $display("%b", po);
# 1  pi=8'b10001000;
#1 $display("%b", po);
# 1  pi=8'b10001001;
#1 $display("%b", po);
# 1  pi=8'b10001010;
#1 $display("%b", po);
# 1  pi=8'b10001011;
#1 $display("%b", po);
# 1  pi=8'b10001100;
#1 $display("%b", po);
# 1  pi=8'b10001101;
#1 $display("%b", po);
# 1  pi=8'b10001110;
#1 $display("%b", po);
# 1  pi=8'b10001111;
#1 $display("%b", po);
# 1  pi=8'b10010000;
#1 $display("%b", po);
# 1  pi=8'b10010001;
#1 $display("%b", po);
# 1  pi=8'b10010010;
#1 $display("%b", po);
# 1  pi=8'b10010011;
#1 $display("%b", po);
# 1  pi=8'b10010100;
#1 $display("%b", po);
# 1  pi=8'b10010101;
#1 $display("%b", po);
# 1  pi=8'b10010110;
#1 $display("%b", po);
# 1  pi=8'b10010111;
#1 $display("%b", po);
# 1  pi=8'b10011000;
#1 $display("%b", po);
# 1  pi=8'b10011001;
#1 $display("%b", po);
# 1  pi=8'b10011010;
#1 $display("%b", po);
# 1  pi=8'b10011011;
#1 $display("%b", po);
# 1  pi=8'b10011100;
#1 $display("%b", po);
# 1  pi=8'b10011101;
#1 $display("%b", po);
# 1  pi=8'b10011110;
#1 $display("%b", po);
# 1  pi=8'b10011111;
#1 $display("%b", po);
# 1  pi=8'b10100000;
#1 $display("%b", po);
# 1  pi=8'b10100001;
#1 $display("%b", po);
# 1  pi=8'b10100010;
#1 $display("%b", po);
# 1  pi=8'b10100011;
#1 $display("%b", po);
# 1  pi=8'b10100100;
#1 $display("%b", po);
# 1  pi=8'b10100101;
#1 $display("%b", po);
# 1  pi=8'b10100110;
#1 $display("%b", po);
# 1  pi=8'b10100111;
#1 $display("%b", po);
# 1  pi=8'b10101000;
#1 $display("%b", po);
# 1  pi=8'b10101001;
#1 $display("%b", po);
# 1  pi=8'b10101010;
#1 $display("%b", po);
# 1  pi=8'b10101011;
#1 $display("%b", po);
# 1  pi=8'b10101100;
#1 $display("%b", po);
# 1  pi=8'b10101101;
#1 $display("%b", po);
# 1  pi=8'b10101110;
#1 $display("%b", po);
# 1  pi=8'b10101111;
#1 $display("%b", po);
# 1  pi=8'b10110000;
#1 $display("%b", po);
# 1  pi=8'b10110001;
#1 $display("%b", po);
# 1  pi=8'b10110010;
#1 $display("%b", po);
# 1  pi=8'b10110011;
#1 $display("%b", po);
# 1  pi=8'b10110100;
#1 $display("%b", po);
# 1  pi=8'b10110101;
#1 $display("%b", po);
# 1  pi=8'b10110110;
#1 $display("%b", po);
# 1  pi=8'b10110111;
#1 $display("%b", po);
# 1  pi=8'b10111000;
#1 $display("%b", po);
# 1  pi=8'b10111001;
#1 $display("%b", po);
# 1  pi=8'b10111010;
#1 $display("%b", po);
# 1  pi=8'b10111011;
#1 $display("%b", po);
# 1  pi=8'b10111100;
#1 $display("%b", po);
# 1  pi=8'b10111101;
#1 $display("%b", po);
# 1  pi=8'b10111110;
#1 $display("%b", po);
# 1  pi=8'b10111111;
#1 $display("%b", po);
# 1  pi=8'b11000000;
#1 $display("%b", po);
# 1  pi=8'b11000001;
#1 $display("%b", po);
# 1  pi=8'b11000010;
#1 $display("%b", po);
# 1  pi=8'b11000011;
#1 $display("%b", po);
# 1  pi=8'b11000100;
#1 $display("%b", po);
# 1  pi=8'b11000101;
#1 $display("%b", po);
# 1  pi=8'b11000110;
#1 $display("%b", po);
# 1  pi=8'b11000111;
#1 $display("%b", po);
# 1  pi=8'b11001000;
#1 $display("%b", po);
# 1  pi=8'b11001001;
#1 $display("%b", po);
# 1  pi=8'b11001010;
#1 $display("%b", po);
# 1  pi=8'b11001011;
#1 $display("%b", po);
# 1  pi=8'b11001100;
#1 $display("%b", po);
# 1  pi=8'b11001101;
#1 $display("%b", po);
# 1  pi=8'b11001110;
#1 $display("%b", po);
# 1  pi=8'b11001111;
#1 $display("%b", po);
# 1  pi=8'b11010000;
#1 $display("%b", po);
# 1  pi=8'b11010001;
#1 $display("%b", po);
# 1  pi=8'b11010010;
#1 $display("%b", po);
# 1  pi=8'b11010011;
#1 $display("%b", po);
# 1  pi=8'b11010100;
#1 $display("%b", po);
# 1  pi=8'b11010101;
#1 $display("%b", po);
# 1  pi=8'b11010110;
#1 $display("%b", po);
# 1  pi=8'b11010111;
#1 $display("%b", po);
# 1  pi=8'b11011000;
#1 $display("%b", po);
# 1  pi=8'b11011001;
#1 $display("%b", po);
# 1  pi=8'b11011010;
#1 $display("%b", po);
# 1  pi=8'b11011011;
#1 $display("%b", po);
# 1  pi=8'b11011100;
#1 $display("%b", po);
# 1  pi=8'b11011101;
#1 $display("%b", po);
# 1  pi=8'b11011110;
#1 $display("%b", po);
# 1  pi=8'b11011111;
#1 $display("%b", po);
# 1  pi=8'b11100000;
#1 $display("%b", po);
# 1  pi=8'b11100001;
#1 $display("%b", po);
# 1  pi=8'b11100010;
#1 $display("%b", po);
# 1  pi=8'b11100011;
#1 $display("%b", po);
# 1  pi=8'b11100100;
#1 $display("%b", po);
# 1  pi=8'b11100101;
#1 $display("%b", po);
# 1  pi=8'b11100110;
#1 $display("%b", po);
# 1  pi=8'b11100111;
#1 $display("%b", po);
# 1  pi=8'b11101000;
#1 $display("%b", po);
# 1  pi=8'b11101001;
#1 $display("%b", po);
# 1  pi=8'b11101010;
#1 $display("%b", po);
# 1  pi=8'b11101011;
#1 $display("%b", po);
# 1  pi=8'b11101100;
#1 $display("%b", po);
# 1  pi=8'b11101101;
#1 $display("%b", po);
# 1  pi=8'b11101110;
#1 $display("%b", po);
# 1  pi=8'b11101111;
#1 $display("%b", po);
# 1  pi=8'b11110000;
#1 $display("%b", po);
# 1  pi=8'b11110001;
#1 $display("%b", po);
# 1  pi=8'b11110010;
#1 $display("%b", po);
# 1  pi=8'b11110011;
#1 $display("%b", po);
# 1  pi=8'b11110100;
#1 $display("%b", po);
# 1  pi=8'b11110101;
#1 $display("%b", po);
# 1  pi=8'b11110110;
#1 $display("%b", po);
# 1  pi=8'b11110111;
#1 $display("%b", po);
# 1  pi=8'b11111000;
#1 $display("%b", po);
# 1  pi=8'b11111001;
#1 $display("%b", po);
# 1  pi=8'b11111010;
#1 $display("%b", po);
# 1  pi=8'b11111011;
#1 $display("%b", po);
# 1  pi=8'b11111100;
#1 $display("%b", po);
# 1  pi=8'b11111101;
#1 $display("%b", po);
# 1  pi=8'b11111110;
#1 $display("%b", po);
end
endmodule
