module mul_i14_o14 (a, b, r);
input [6:0] a, b;
output [13:0] r;


assign r = a * b;

endmodule 
