// Benchmark "circuit" written by ABC on Mon Apr 25 13:08:35 2022

module circuit ( 
    g0, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15,
    g963, g962, g961, g960, g959, g958, g957, g956, g955, g954, g953, g952,
    g951, g950, g949, g948, g947, g946  );
  input  g0, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14,
    g15;
  output g963, g962, g961, g960, g959, g958, g957, g956, g955, g954, g953,
    g952, g951, g950, g949, g948, g947, g946;
  wire g16, g17, g18, g19, g20, g21, g22, g23, g24, g25, g26, g27, g28, g29,
    g30, g31, g32, g33, g34, g35, g36, g37, g38, g39, g40, g41, g42, g43,
    g44, g45, g46, g47, g48, g49, g50, g51, g52, g53, g54, g55, g56, g57,
    g58, g59, g60, g61, g62, g63, g64, g65, g66, g67, g68, g69, g70, g71,
    g72, g73, g74, g75, g76, g77, g78, g79, g80, g81, g82, g83, g84, g85,
    g86, g87, g88, g89, g90, g91, g92, g93, g94, g95, g96, g97, g98, g99,
    g100, g101, g102, g103, g104, g105, g106, g107, g108, g109, g110, g111,
    g112, g113, g114, g115, g116, g117, g118, g119, g120, g121, g122, g123,
    g124, g125, g126, g127, g128, g129, g130, g131, g132, g133, g134, g135,
    g136, g137, g138, g139, g140, g141, g142, g143, g144, g145, g146, g147,
    g148, g149, g150, g151, g152, g153, g154, g155, g156, g157, g158, g159,
    g160, g161, g162, g163, g164, g165, g166, g167, g168, g169, g170, g171,
    g172, g173, g174, g175, g176, g177, g178, g179, g180, g181, g182, g183,
    g184, g185, g186, g187, g188, g189, g190, g191, g192, g193, g194, g195,
    g196, g197, g198, g199, g200, g201, g202, g203, g204, g205, g206, g207,
    g208, g209, g210, g211, g212, g213, g214, g215, g216, g217, g218, g219,
    g220, g221, g222, g223, g224, g225, g226, g227, g228, g229, g230, g231,
    g232, g233, g234, g235, g236, g237, g238, g239, g240, g241, g242, g243,
    g244, g245, g246, g247, g248, g249, g250, g251, g252, g253, g254, g255,
    g256, g257, g258, g259, g260, g261, g262, g263, g264, g265, g266, g267,
    g268, g269, g270, g271, g272, g273, g274, g275, g276, g277, g278, g279,
    g280, g281, g282, g283, g284, g285, g286, g287, g288, g289, g290, g291,
    g292, g293, g294, g295, g296, g297, g298, g299, g300, g301, g302, g303,
    g304, g305, g306, g307, g308, g309, g310, g311, g312, g313, g314, g315,
    g316, g317, g318, g319, g320, g321, g322, g323, g324, g325, g326, g327,
    g328, g329, g330, g331, g332, g333, g334, g335, g336, g337, g338, g339,
    g340, g341, g342, g343, g344, g345, g346, g347, g348, g349, g350, g351,
    g352, g353, g354, g355, g356, g357, g358, g359, g360, g361, g362, g363,
    g364, g365, g366, g367, g368, g369, g370, g371, g372, g373, g374, g375,
    g376, g377, g378, g379, g380, g381, g382, g383, g384, g385, g386, g387,
    g388, g389, g390, g391, g392, g393, g394, g395, g396, g397, g398, g399,
    g400, g401, g402, g403, g404, g405, g406, g407, g408, g409, g410, g411,
    g412, g413, g414, g415, g416, g417, g418, g419, g420, g421, g422, g423,
    g424, g425, g426, g427, g428, g429, g430, g431, g432, g433, g434, g435,
    g436, g437, g438, g439, g440, g441, g442, g443, g444, g445, g446, g447,
    g448, g449, g450, g451, g452, g453, g454, g455, g456, g457, g458, g459,
    g460, g461, g462, g463, g464, g465, g466, g467, g468, g469, g470, g471,
    g472, g473, g474, g475, g476, g477, g478, g479, g480, g481, g482, g483,
    g484, g485, g486, g487, g488, g489, g490, g491, g492, g493, g494, g495,
    g496, g497, g498, g499, g500, g501, g502, g503, g504, g505, g506, g507,
    g508, g509, g510, g511, g512, g513, g514, g515, g516, g517, g518, g519,
    g520, g521, g522, g523, g524, g525, g526, g527, g528, g529, g530, g531,
    g532, g533, g534, g535, g536, g537, g538, g539, g540, g541, g542, g543,
    g544, g545, g546, g547, g548, g549, g550, g551, g552, g553, g554, g555,
    g556, g557, g558, g559, g560, g561, g562, g563, g564, g565, g566, g567,
    g568, g569, g570, g571, g572, g573, g574, g575, g576, g577, g578, g579,
    g580, g581, g582, g583, g584, g585, g586, g587, g588, g589, g590, g591,
    g592, g593, g594, g595, g596, g597, g598, g599, g600, g601, g602, g603,
    g604, g605, g606, g607, g608, g609, g610, g611, g612, g613, g614, g615,
    g616, g617, g618, g619, g620, g621, g622, g623, g624, g625, g626, g627,
    g628, g629, g630, g631, g632, g633, g634, g635, g636, g637, g638, g639,
    g640, g641, g642, g643, g644, g645, g646, g647, g648, g649, g650, g651,
    g652, g653, g654, g655, g656, g657, g658, g659, g660, g661, g662, g663,
    g664, g665, g666, g667, g668, g669, g670, g671, g672, g673, g674, g675,
    g676, g677, g678, g679, g680, g681, g682, g683, g684, g685, g686, g687,
    g688, g689, g690, g691, g692, g693, g694, g695, g696, g697, g698, g699,
    g700, g701, g702, g703, g704, g705, g706, g707, g708, g709, g710, g711,
    g712, g713, g714, g715, g716, g717, g718, g719, g720, g721, g722, g723,
    g724, g725, g726, g727, g728, g729, g730, g731, g732, g733, g734, g735,
    g736, g737, g738, g739, g740, g741, g742, g743, g744, g745, g746, g747,
    g748, g749, g750, g751, g752, g753, g754, g755, g756, g757, g758, g759,
    g760, g761, g762, g763, g764, g765, g766, g767, g768, g769, g770, g771,
    g772, g773, g774, g775, g776, g777, g778, g779, g780, g781, g782, g783,
    g784, g785, g786, g787, g788, g789, g790, g791, g792, g793, g794, g795,
    g796, g797, g798, g799, g800, g801, g802, g803, g804, g805, g806, g807,
    g808, g809, g810, g811, g812, g813, g814, g815, g816, g817, g818, g819,
    g820, g821, g822, g823, g824, g825, g826, g827, g828, g829, g830, g831,
    g832, g833, g834, g835, g836, g837, g838, g839, g840, g841, g842, g843,
    g844, g845, g846, g847, g848, g849, g850, g851, g852, g853, g854, g855,
    g856, g857, g858, g859, g860, g861, g862, g863, g864, g865, g866, g867,
    g868, g869, g870, g871, g872, g873, g874, g875, g876, g877, g878, g879,
    g880, g881, g882, g883, g884, g885, g886, g887, g888, g889, g890, g891,
    g892, g893, g894, g895, g896, g897, g898, g899, g900, g901, g902, g903,
    g904, g905, g906, g907, g908, g909, g910, g911, g912, g913, g914, g915,
    g916, g917, g918, g919, g920, g921, g922, g923, g924, g925, g926, g927,
    g928, g929, g930, g931, g932, g933, g934, g935, g936, g937, g938, g939,
    g940, g941, g942, g943, g944, g945;
  assign g16 = ~g15;
  assign g17 = ~g14;
  assign g18 = ~g13;
  assign g19 = ~g12;
  assign g20 = ~g11;
  assign g21 = ~g10;
  assign g22 = ~g9;
  assign g23 = ~g8;
  assign g24 = ~g7;
  assign g25 = ~g15 | ~g24;
  assign g26 = ~g7 | ~g16;
  assign g27 = ~g25 | ~g26;
  assign g28 = ~g27;
  assign g29 = ~g6;
  assign g30 = ~g14 | ~g29;
  assign g31 = ~g6 | ~g17;
  assign g32 = ~g30 | ~g31;
  assign g33 = ~g32;
  assign g34 = ~g5;
  assign g35 = ~g13 | ~g34;
  assign g36 = ~g5 | ~g18;
  assign g37 = ~g35 | ~g36;
  assign g38 = ~g37;
  assign g39 = ~g4;
  assign g40 = ~g12 | ~g39;
  assign g41 = ~g4 | ~g19;
  assign g42 = ~g40 | ~g41;
  assign g43 = ~g42;
  assign g44 = ~g3;
  assign g45 = ~g11 | ~g44;
  assign g46 = ~g3 | ~g20;
  assign g47 = ~g45 | ~g46;
  assign g48 = ~g47;
  assign g49 = ~g2;
  assign g50 = ~g10 | ~g49;
  assign g51 = ~g2 | ~g21;
  assign g52 = ~g50 | ~g51;
  assign g53 = ~g52;
  assign g54 = ~g1;
  assign g55 = ~g9 | ~g54;
  assign g56 = ~g1 | ~g22;
  assign g57 = ~g55 | ~g56;
  assign g58 = ~g57;
  assign g59 = ~g0 | ~g23;
  assign g60 = ~g0 & ~g23;
  assign g61 = ~g54 | ~g60;
  assign g62 = ~g22 | ~g61;
  assign g63 = ~g58 | ~g60;
  assign g64 = ~g60;
  assign g65 = ~g1 | ~g64;
  assign g66 = ~g62 | ~g65;
  assign g67 = ~g2 | ~g66;
  assign g68 = ~g66;
  assign g69 = ~g49 | ~g68;
  assign g70 = ~g21 | ~g69;
  assign g71 = ~g67 | ~g70;
  assign g72 = ~g3 | ~g71;
  assign g73 = ~g71;
  assign g74 = ~g44 | ~g73;
  assign g75 = ~g20 | ~g74;
  assign g76 = ~g72 | ~g75;
  assign g77 = ~g4 | ~g76;
  assign g78 = ~g76;
  assign g79 = ~g39 | ~g78;
  assign g80 = ~g19 | ~g79;
  assign g81 = ~g77 | ~g80;
  assign g82 = ~g5 | ~g81;
  assign g83 = ~g81;
  assign g84 = ~g34 | ~g83;
  assign g85 = ~g18 | ~g84;
  assign g86 = ~g82 | ~g85;
  assign g87 = ~g6 | ~g86;
  assign g88 = ~g86;
  assign g89 = ~g29 | ~g88;
  assign g90 = ~g17 | ~g89;
  assign g91 = ~g87 | ~g90;
  assign g92 = ~g7 | ~g91;
  assign g93 = ~g91;
  assign g94 = ~g24 | ~g93;
  assign g95 = ~g16 | ~g94;
  assign g96 = ~g92 | ~g95;
  assign g97 = ~g96;
  assign g98 = ~g28 | ~g97;
  assign g99 = ~g27 | ~g96;
  assign g100 = ~g98 | ~g99;
  assign g101 = ~g100 | ~g100;
  assign g102 = ~g101;
  assign g103 = ~g28 | ~g93;
  assign g104 = ~g27 | ~g91;
  assign g105 = ~g103 | ~g104;
  assign g106 = ~g100 | ~g105;
  assign g107 = ~g106;
  assign g108 = 1'b0;
  assign g109 = ~g100 | ~g105;
  assign g110 = ~g106 | ~g109;
  assign g111 = ~g105 | ~g105;
  assign g112 = ~g111;
  assign g113 = ~g33 | ~g88;
  assign g114 = ~g32 | ~g86;
  assign g115 = ~g113 | ~g114;
  assign g116 = ~g100 | ~g115;
  assign g117 = ~g116;
  assign g118 = ~g111 | ~g117;
  assign g119 = ~g100 | ~g115;
  assign g120 = ~g112 | ~g119;
  assign g121 = ~g118 | ~g120;
  assign g122 = ~g121;
  assign g123 = ~g116 | ~g122;
  assign g124 = ~g120 | ~g123;
  assign g125 = ~g108 & ~g124;
  assign g126 = ~g125;
  assign g127 = ~g108 | ~g124;
  assign g128 = ~g110 | ~g127;
  assign g129 = ~g102 | ~g128;
  assign g130 = 1'b0;
  assign g131 = ~g101 | ~g130;
  assign g132 = ~g129 | ~g131;
  assign g133 = ~g132;
  assign g134 = ~g126 | ~g127;
  assign g135 = ~g134;
  assign g136 = ~g117 | ~g122;
  assign g137 = ~g116 | ~g121;
  assign g138 = ~g136 | ~g137;
  assign g139 = ~g105 | ~g115;
  assign g140 = ~g139;
  assign g141 = ~g105 | ~g115;
  assign g142 = ~g115 | ~g115;
  assign g143 = ~g142;
  assign g144 = ~g38 | ~g83;
  assign g145 = ~g37 | ~g81;
  assign g146 = ~g144 | ~g145;
  assign g147 = ~g100 | ~g146;
  assign g148 = ~g147;
  assign g149 = ~g139 | ~g148;
  assign g150 = ~g100 | ~g146;
  assign g151 = ~g140 | ~g150;
  assign g152 = ~g149 | ~g151;
  assign g153 = ~g152;
  assign g154 = ~g147 | ~g153;
  assign g155 = ~g151 | ~g154;
  assign g156 = ~g138 & ~g155;
  assign g157 = ~g156;
  assign g158 = ~g138 | ~g155;
  assign g159 = ~g157 | ~g158;
  assign g160 = ~g159;
  assign g161 = ~g148 | ~g153;
  assign g162 = ~g147 | ~g152;
  assign g163 = ~g161 | ~g162;
  assign g164 = ~g163;
  assign g165 = ~g105 | ~g146;
  assign g166 = ~g165;
  assign g167 = 1'b0;
  assign g168 = ~g115 | ~g146;
  assign g169 = ~g115 | ~g146;
  assign g170 = ~g169;
  assign g171 = ~g146 | ~g146;
  assign g172 = ~g171;
  assign g173 = ~g43 | ~g78;
  assign g174 = ~g42 | ~g76;
  assign g175 = ~g173 | ~g174;
  assign g176 = ~g100 | ~g175;
  assign g177 = ~g176;
  assign g178 = ~g142 | ~g177;
  assign g179 = ~g100 | ~g175;
  assign g180 = ~g143 | ~g179;
  assign g181 = ~g178 | ~g180;
  assign g182 = ~g181;
  assign g183 = ~g176 | ~g182;
  assign g184 = ~g180 | ~g183;
  assign g185 = ~g140 | ~g184;
  assign g186 = ~g184;
  assign g187 = ~g141 | ~g186;
  assign g188 = ~g185 | ~g187;
  assign g189 = ~g188;
  assign g190 = ~g177 | ~g182;
  assign g191 = ~g176 | ~g181;
  assign g192 = ~g190 | ~g191;
  assign g193 = ~g192;
  assign g194 = ~g105 | ~g175;
  assign g195 = ~g194;
  assign g196 = ~g170 | ~g195;
  assign g197 = ~g169 | ~g195;
  assign g198 = ~g105 | ~g175;
  assign g199 = ~g170 | ~g198;
  assign g200 = ~g197 | ~g199;
  assign g201 = ~g195 | ~g200;
  assign g202 = ~g196 | ~g201;
  assign g203 = ~g167 & ~g202;
  assign g204 = ~g203;
  assign g205 = ~g167 | ~g202;
  assign g206 = ~g165 | ~g205;
  assign g207 = ~g189 | ~g206;
  assign g208 = ~g185 | ~g207;
  assign g209 = ~g160 | ~g208;
  assign g210 = ~g158 | ~g209;
  assign g211 = ~g135 | ~g210;
  assign g212 = ~g210;
  assign g213 = ~g135 | ~g212;
  assign g214 = ~g134 | ~g210;
  assign g215 = ~g213 | ~g214;
  assign g216 = ~g208;
  assign g217 = ~g160 | ~g216;
  assign g218 = ~g159 | ~g208;
  assign g219 = ~g217 | ~g218;
  assign g220 = ~g206;
  assign g221 = ~g189 | ~g220;
  assign g222 = ~g188 | ~g206;
  assign g223 = ~g221 | ~g222;
  assign g224 = ~g163 | ~g223;
  assign g225 = ~g223;
  assign g226 = ~g163 | ~g225;
  assign g227 = ~g164 | ~g223;
  assign g228 = ~g226 | ~g227;
  assign g229 = ~g204 | ~g205;
  assign g230 = ~g229;
  assign g231 = ~g200;
  assign g232 = ~g195 | ~g231;
  assign g233 = ~g194 | ~g200;
  assign g234 = ~g232 | ~g233;
  assign g235 = ~g115 | ~g175;
  assign g236 = ~g235;
  assign g237 = ~g146 | ~g175;
  assign g238 = ~g237;
  assign g239 = ~g175 | ~g175;
  assign g240 = ~g239;
  assign g241 = ~g146 | ~g175;
  assign g242 = ~g241;
  assign g243 = ~g115 | ~g175;
  assign g244 = ~g48 | ~g73;
  assign g245 = ~g47 | ~g71;
  assign g246 = ~g244 | ~g245;
  assign g247 = ~g100 | ~g246;
  assign g248 = ~g247;
  assign g249 = ~g168 | ~g248;
  assign g250 = ~g100 | ~g246;
  assign g251 = ~g170 | ~g250;
  assign g252 = ~g249 | ~g251;
  assign g253 = ~g252;
  assign g254 = ~g247 | ~g253;
  assign g255 = ~g251 | ~g254;
  assign g256 = ~g230 | ~g255;
  assign g257 = ~g255;
  assign g258 = ~g230 | ~g257;
  assign g259 = ~g229 | ~g255;
  assign g260 = ~g258 | ~g259;
  assign g261 = ~g192 | ~g260;
  assign g262 = ~g256 | ~g261;
  assign g263 = ~g228 & ~g262;
  assign g264 = ~g263;
  assign g265 = ~g228 | ~g262;
  assign g266 = ~g224 | ~g265;
  assign g267 = ~g219 & ~g266;
  assign g268 = ~g267;
  assign g269 = ~g219 | ~g266;
  assign g270 = ~g268 | ~g269;
  assign g271 = ~g270;
  assign g272 = ~g264 | ~g265;
  assign g273 = ~g272;
  assign g274 = ~g260;
  assign g275 = ~g192 | ~g274;
  assign g276 = ~g193 | ~g260;
  assign g277 = ~g275 | ~g276;
  assign g278 = ~g277;
  assign g279 = ~g248 | ~g253;
  assign g280 = ~g247 | ~g252;
  assign g281 = ~g279 | ~g280;
  assign g282 = ~g281;
  assign g283 = ~g246 | ~g246;
  assign g284 = ~g283;
  assign g285 = ~g105 | ~g246;
  assign g286 = ~g236 | ~g285;
  assign g287 = ~g285;
  assign g288 = ~g236 | ~g287;
  assign g289 = ~g235 | ~g287;
  assign g290 = ~g286 | ~g289;
  assign g291 = ~g175 | ~g246;
  assign g292 = ~g291;
  assign g293 = 1'b0;
  assign g294 = ~g115 | ~g246;
  assign g295 = ~g294;
  assign g296 = ~g146 | ~g246;
  assign g297 = ~g296;
  assign g298 = ~g146 | ~g246;
  assign g299 = ~g105 | ~g246;
  assign g300 = ~g53 | ~g68;
  assign g301 = ~g52 | ~g66;
  assign g302 = ~g300 | ~g301;
  assign g303 = ~g302 | ~g302;
  assign g304 = ~g303;
  assign g305 = ~g246 | ~g302;
  assign g306 = ~g246 | ~g302;
  assign g307 = ~g306;
  assign g308 = ~g146 | ~g302;
  assign g309 = ~g146 | ~g302;
  assign g310 = ~g309;
  assign g311 = ~g100 | ~g302;
  assign g312 = ~g311;
  assign g313 = ~g243 | ~g312;
  assign g314 = ~g175 | ~g302;
  assign g315 = ~g314;
  assign g316 = ~g175 | ~g302;
  assign g317 = ~g316;
  assign g318 = ~g105 | ~g302;
  assign g319 = ~g237 | ~g318;
  assign g320 = ~g172 | ~g319;
  assign g321 = ~g319;
  assign g322 = ~g171 | ~g321;
  assign g323 = ~g320 | ~g322;
  assign g324 = ~g323;
  assign g325 = ~g311 | ~g324;
  assign g326 = ~g320 | ~g325;
  assign g327 = ~g326;
  assign g328 = ~g312 | ~g324;
  assign g329 = ~g311 | ~g323;
  assign g330 = ~g328 | ~g329;
  assign g331 = ~g330;
  assign g332 = ~g238 | ~g318;
  assign g333 = ~g115 | ~g302;
  assign g334 = ~g333;
  assign g335 = ~g297 | ~g334;
  assign g336 = ~g115 | ~g335;
  assign g337 = ~g336;
  assign g338 = ~g246 | ~g337;
  assign g339 = ~g298 | ~g334;
  assign g340 = ~g297 | ~g333;
  assign g341 = ~g339 | ~g340;
  assign g342 = ~g297 | ~g341;
  assign g343 = ~g341;
  assign g344 = ~g297 | ~g343;
  assign g345 = ~g296 | ~g341;
  assign g346 = ~g344 | ~g345;
  assign g347 = ~g346;
  assign g348 = ~g115 | ~g302;
  assign g349 = ~g105 | ~g302;
  assign g350 = ~g349;
  assign g351 = ~g237 | ~g350;
  assign g352 = ~g332 | ~g351;
  assign g353 = ~g338 & ~g352;
  assign g354 = ~g353;
  assign g355 = ~g335 | ~g354;
  assign g356 = ~g355;
  assign g357 = ~g338 | ~g352;
  assign g358 = ~g354 | ~g357;
  assign g359 = ~g358;
  assign g360 = ~g242 | ~g350;
  assign g361 = ~g241 | ~g350;
  assign g362 = ~g242 | ~g349;
  assign g363 = ~g361 | ~g362;
  assign g364 = ~g100 | ~g302;
  assign g365 = ~g236 | ~g364;
  assign g366 = ~g313 | ~g365;
  assign g367 = ~g366;
  assign g368 = ~g287 | ~g367;
  assign g369 = ~g365 | ~g368;
  assign g370 = ~g326 | ~g369;
  assign g371 = ~g369;
  assign g372 = ~g326 | ~g371;
  assign g373 = ~g327 | ~g369;
  assign g374 = ~g372 | ~g373;
  assign g375 = ~g299 | ~g366;
  assign g376 = ~g368 | ~g375;
  assign g377 = ~g376;
  assign g378 = ~g57 | ~g64;
  assign g379 = ~g63 | ~g378;
  assign g380 = ~g302 | ~g379;
  assign g381 = ~g302 | ~g379;
  assign g382 = ~g381;
  assign g383 = ~g379 | ~g379;
  assign g384 = ~g383;
  assign g385 = ~g246 | ~g379;
  assign g386 = ~g385;
  assign g387 = ~g304 | ~g386;
  assign g388 = ~g303 | ~g386;
  assign g389 = ~g304 | ~g385;
  assign g390 = ~g388 | ~g389;
  assign g391 = ~g246 | ~g379;
  assign g392 = ~g175 | ~g379;
  assign g393 = ~g392;
  assign g394 = ~g307 | ~g393;
  assign g395 = ~g305 | ~g393;
  assign g396 = ~g175 | ~g379;
  assign g397 = ~g307 | ~g396;
  assign g398 = ~g395 | ~g397;
  assign g399 = ~g398;
  assign g400 = ~g307 | ~g399;
  assign g401 = ~g306 | ~g398;
  assign g402 = ~g400 | ~g401;
  assign g403 = ~g307 | ~g398;
  assign g404 = ~g394 | ~g403;
  assign g405 = ~g284 | ~g404;
  assign g406 = ~g404;
  assign g407 = ~g283 | ~g406;
  assign g408 = ~g405 | ~g407;
  assign g409 = ~g408;
  assign g410 = ~g115 | ~g379;
  assign g411 = ~g410;
  assign g412 = ~g310 | ~g411;
  assign g413 = ~g308 | ~g411;
  assign g414 = ~g310 | ~g410;
  assign g415 = ~g413 | ~g414;
  assign g416 = ~g415;
  assign g417 = ~g310 | ~g416;
  assign g418 = ~g309 | ~g415;
  assign g419 = ~g417 | ~g418;
  assign g420 = 1'b0;
  assign g421 = ~g310 | ~g415;
  assign g422 = ~g412 | ~g421;
  assign g423 = ~g422;
  assign g424 = ~g146 | ~g379;
  assign g425 = ~g424;
  assign g426 = ~g146 | ~g379;
  assign g427 = ~g426;
  assign g428 = ~g315 | ~g427;
  assign g429 = ~g314 | ~g427;
  assign g430 = ~g315 | ~g426;
  assign g431 = ~g429 | ~g430;
  assign g432 = ~g431;
  assign g433 = ~g317 | ~g432;
  assign g434 = ~g316 | ~g431;
  assign g435 = ~g433 | ~g434;
  assign g436 = ~g435;
  assign g437 = ~g408 | ~g436;
  assign g438 = ~g409 | ~g435;
  assign g439 = ~g437 | ~g438;
  assign g440 = ~g439;
  assign g441 = ~g405 | ~g438;
  assign g442 = ~g317 | ~g431;
  assign g443 = ~g428 | ~g442;
  assign g444 = ~g293 & ~g443;
  assign g445 = ~g444;
  assign g446 = ~g293 | ~g443;
  assign g447 = ~g291 | ~g446;
  assign g448 = ~g445 | ~g446;
  assign g449 = ~g448;
  assign g450 = ~g100 | ~g379;
  assign g451 = ~g450;
  assign g452 = ~g294 | ~g451;
  assign g453 = ~g100 | ~g379;
  assign g454 = ~g295 | ~g453;
  assign g455 = ~g452 | ~g454;
  assign g456 = ~g455;
  assign g457 = ~g450 | ~g456;
  assign g458 = ~g454 | ~g457;
  assign g459 = ~g290 & ~g458;
  assign g460 = ~g459;
  assign g461 = ~g290 | ~g458;
  assign g462 = ~g288 | ~g461;
  assign g463 = ~g234 & ~g462;
  assign g464 = ~g463;
  assign g465 = ~g234 | ~g462;
  assign g466 = ~g464 | ~g465;
  assign g467 = ~g466;
  assign g468 = ~g281 | ~g467;
  assign g469 = ~g465 | ~g468;
  assign g470 = ~g469;
  assign g471 = ~g282 | ~g466;
  assign g472 = ~g468 | ~g471;
  assign g473 = ~g472;
  assign g474 = ~g460 | ~g461;
  assign g475 = ~g474;
  assign g476 = ~g355 | ~g475;
  assign g477 = ~g356 | ~g475;
  assign g478 = ~g355 | ~g474;
  assign g479 = ~g477 | ~g478;
  assign g480 = ~g330 | ~g479;
  assign g481 = ~g476 | ~g480;
  assign g482 = ~g374 & ~g481;
  assign g483 = ~g482;
  assign g484 = ~g374 | ~g481;
  assign g485 = ~g370 | ~g484;
  assign g486 = ~g469 | ~g485;
  assign g487 = ~g470 | ~g485;
  assign g488 = ~g485;
  assign g489 = ~g469 | ~g488;
  assign g490 = ~g487 | ~g489;
  assign g491 = ~g277 | ~g490;
  assign g492 = ~g486 | ~g491;
  assign g493 = ~g273 | ~g492;
  assign g494 = ~g492;
  assign g495 = ~g273 | ~g494;
  assign g496 = ~g272 | ~g492;
  assign g497 = ~g495 | ~g496;
  assign g498 = ~g490;
  assign g499 = ~g277 | ~g498;
  assign g500 = ~g278 | ~g490;
  assign g501 = ~g499 | ~g500;
  assign g502 = ~g483 | ~g484;
  assign g503 = ~g473 | ~g502;
  assign g504 = ~g502;
  assign g505 = ~g473 | ~g504;
  assign g506 = ~g472 | ~g504;
  assign g507 = ~g503 | ~g506;
  assign g508 = ~g479;
  assign g509 = ~g330 | ~g508;
  assign g510 = ~g331 | ~g479;
  assign g511 = ~g509 | ~g510;
  assign g512 = ~g511;
  assign g513 = ~g451 | ~g456;
  assign g514 = ~g450 | ~g455;
  assign g515 = ~g513 | ~g514;
  assign g516 = ~g359 | ~g515;
  assign g517 = ~g515;
  assign g518 = ~g358 | ~g517;
  assign g519 = ~g516 | ~g518;
  assign g520 = ~g519;
  assign g521 = ~g115 | ~g379;
  assign g522 = ~g105 | ~g379;
  assign g523 = ~g522;
  assign g524 = 1'b0;
  assign g525 = ~g524;
  assign g526 = ~g240 | ~g525;
  assign g527 = ~g239 | ~g524;
  assign g528 = ~g526 | ~g527;
  assign g529 = ~g528;
  assign g530 = ~g240 | ~g524;
  assign g531 = ~g522 | ~g530;
  assign g532 = ~g363 & ~g531;
  assign g533 = ~g532;
  assign g534 = ~g363 | ~g531;
  assign g535 = ~g533 | ~g534;
  assign g536 = ~g535;
  assign g537 = ~g360 | ~g534;
  assign g538 = ~g377 | ~g537;
  assign g539 = ~g537;
  assign g540 = ~g377 | ~g539;
  assign g541 = ~g376 | ~g537;
  assign g542 = ~g540 | ~g541;
  assign g543 = ~g59 | ~g64;
  assign g544 = ~g302 | ~g543;
  assign g545 = ~g544;
  assign g546 = ~g383 | ~g545;
  assign g547 = ~g384 | ~g545;
  assign g548 = ~g379 | ~g543;
  assign g549 = ~g548;
  assign g550 = 1'b0;
  assign g551 = ~g549 | ~g549;
  assign g552 = ~g551;
  assign g553 = ~g175 | ~g543;
  assign g554 = ~g246 | ~g543;
  assign g555 = ~g382 | ~g554;
  assign g556 = ~g554;
  assign g557 = ~g380 | ~g556;
  assign g558 = ~g555 | ~g557;
  assign g559 = ~g558;
  assign g560 = ~g381 | ~g556;
  assign g561 = ~g382 | ~g556;
  assign g562 = ~g561;
  assign g563 = ~g382 | ~g556;
  assign g564 = ~g547 | ~g563;
  assign g565 = ~g390 & ~g564;
  assign g566 = ~g565;
  assign g567 = ~g390 | ~g564;
  assign g568 = ~g566 | ~g567;
  assign g569 = ~g568;
  assign g570 = ~g387 | ~g567;
  assign g571 = ~g402 & ~g570;
  assign g572 = ~g571;
  assign g573 = ~g402 | ~g570;
  assign g574 = ~g572 | ~g573;
  assign g575 = ~g574;
  assign g576 = ~g246 | ~g543;
  assign g577 = ~g382 | ~g576;
  assign g578 = ~g560 | ~g577;
  assign g579 = ~g547 & ~g578;
  assign g580 = ~g579;
  assign g581 = ~g547 | ~g578;
  assign g582 = ~g580 | ~g581;
  assign g583 = ~g558 | ~g582;
  assign g584 = ~g582;
  assign g585 = ~g558 | ~g584;
  assign g586 = ~g559 | ~g582;
  assign g587 = ~g585 | ~g586;
  assign g588 = ~g302 | ~g543;
  assign g589 = ~g384 | ~g588;
  assign g590 = ~g546 | ~g589;
  assign g591 = ~g545 | ~g590;
  assign g592 = ~g590;
  assign g593 = 1'b0;
  assign g594 = 1'b0;
  assign g595 = ~g593 | ~g594;
  assign g596 = 1'b0;
  assign g597 = 1'b0;
  assign g598 = 1'b0;
  assign g599 = 1'b0;
  assign g600 = ~g552 | ~g595;
  assign g601 = ~g591 | ~g600;
  assign g602 = ~g587 & ~g601;
  assign g603 = ~g587 | ~g601;
  assign g604 = ~g603;
  assign g605 = ~g602 & ~g604;
  assign g606 = ~g583 | ~g603;
  assign g607 = ~g606;
  assign g608 = ~g146 | ~g543;
  assign g609 = ~g608;
  assign g610 = ~g392 | ~g609;
  assign g611 = ~g393 | ~g609;
  assign g612 = ~g611;
  assign g613 = ~g175 | ~g543;
  assign g614 = ~g386 | ~g613;
  assign g615 = ~g613;
  assign g616 = ~g391 | ~g615;
  assign g617 = ~g614 | ~g616;
  assign g618 = ~g615 | ~g617;
  assign g619 = ~g617;
  assign g620 = ~g615 | ~g619;
  assign g621 = ~g553 | ~g617;
  assign g622 = ~g620 | ~g621;
  assign g623 = 1'b0;
  assign g624 = ~g562 | ~g623;
  assign g625 = ~g561 | ~g622;
  assign g626 = ~g624 | ~g625;
  assign g627 = ~g569 | ~g626;
  assign g628 = ~g626;
  assign g629 = ~g568 | ~g628;
  assign g630 = ~g627 | ~g629;
  assign g631 = ~g606 | ~g630;
  assign g632 = ~g630;
  assign g633 = ~g607 | ~g632;
  assign g634 = ~g631 | ~g633;
  assign g635 = ~g606 | ~g632;
  assign g636 = ~g627 | ~g635;
  assign g637 = ~g562 | ~g622;
  assign g638 = ~g618 | ~g637;
  assign g639 = ~g638;
  assign g640 = ~g575 | ~g639;
  assign g641 = ~g574 | ~g638;
  assign g642 = ~g640 | ~g641;
  assign g643 = ~g642;
  assign g644 = ~g575 | ~g638;
  assign g645 = ~g573 | ~g644;
  assign g646 = ~g386 | ~g615;
  assign g647 = ~g646;
  assign g648 = ~g115 | ~g543;
  assign g649 = ~g648;
  assign g650 = ~g146 | ~g543;
  assign g651 = ~g393 | ~g650;
  assign g652 = ~g610 | ~g651;
  assign g653 = ~g609 | ~g652;
  assign g654 = ~g652;
  assign g655 = ~g609 | ~g654;
  assign g656 = ~g608 | ~g652;
  assign g657 = ~g655 | ~g656;
  assign g658 = 1'b0;
  assign g659 = ~g647 | ~g658;
  assign g660 = ~g646 | ~g657;
  assign g661 = ~g659 | ~g660;
  assign g662 = ~g642 | ~g661;
  assign g663 = ~g643 | ~g661;
  assign g664 = ~g661;
  assign g665 = ~g642 | ~g664;
  assign g666 = ~g663 | ~g665;
  assign g667 = ~g636 & ~g666;
  assign g668 = ~g636 | ~g666;
  assign g669 = ~g668;
  assign g670 = ~g667 & ~g669;
  assign g671 = ~g662 | ~g668;
  assign g672 = ~g671;
  assign g673 = ~g647 | ~g657;
  assign g674 = ~g653 | ~g673;
  assign g675 = ~g440 | ~g674;
  assign g676 = ~g674;
  assign g677 = ~g440 | ~g676;
  assign g678 = ~g439 | ~g674;
  assign g679 = ~g677 | ~g678;
  assign g680 = ~g679;
  assign g681 = ~g105 | ~g543;
  assign g682 = ~g681;
  assign g683 = ~g521 | ~g682;
  assign g684 = ~g411 | ~g682;
  assign g685 = ~g346 | ~g684;
  assign g686 = ~g684;
  assign g687 = ~g347 | ~g686;
  assign g688 = ~g685 | ~g687;
  assign g689 = ~g688;
  assign g690 = ~g346 | ~g686;
  assign g691 = ~g342 | ~g690;
  assign g692 = ~g115 | ~g543;
  assign g693 = ~g425 | ~g692;
  assign g694 = ~g692;
  assign g695 = ~g424 | ~g694;
  assign g696 = ~g693 | ~g695;
  assign g697 = ~g649 | ~g696;
  assign g698 = ~g696;
  assign g699 = ~g649 | ~g698;
  assign g700 = ~g648 | ~g696;
  assign g701 = ~g699 | ~g700;
  assign g702 = 1'b0;
  assign g703 = ~g612 | ~g702;
  assign g704 = ~g611 | ~g701;
  assign g705 = ~g703 | ~g704;
  assign g706 = ~g680 | ~g705;
  assign g707 = ~g705;
  assign g708 = ~g679 | ~g707;
  assign g709 = ~g706 | ~g708;
  assign g710 = ~g645 & ~g709;
  assign g711 = ~g710;
  assign g712 = ~g645 | ~g709;
  assign g713 = ~g711 | ~g712;
  assign g714 = ~g671 | ~g713;
  assign g715 = ~g713;
  assign g716 = ~g672 | ~g715;
  assign g717 = ~g714 | ~g716;
  assign g718 = ~g671 | ~g715;
  assign g719 = ~g712 | ~g718;
  assign g720 = ~g679 | ~g705;
  assign g721 = ~g675 | ~g720;
  assign g722 = ~g721;
  assign g723 = ~g612 | ~g701;
  assign g724 = ~g697 | ~g723;
  assign g725 = ~g449 | ~g724;
  assign g726 = ~g724;
  assign g727 = ~g449 | ~g726;
  assign g728 = ~g448 | ~g724;
  assign g729 = ~g727 | ~g728;
  assign g730 = ~g729;
  assign g731 = ~g425 | ~g694;
  assign g732 = ~g731;
  assign g733 = ~g105 | ~g543;
  assign g734 = ~g411 | ~g733;
  assign g735 = ~g683 | ~g734;
  assign g736 = ~g682 | ~g735;
  assign g737 = ~g735;
  assign g738 = ~g682 | ~g737;
  assign g739 = ~g681 | ~g735;
  assign g740 = ~g738 | ~g739;
  assign g741 = 1'b0;
  assign g742 = ~g732 | ~g741;
  assign g743 = ~g731 | ~g740;
  assign g744 = ~g742 | ~g743;
  assign g745 = ~g419 | ~g744;
  assign g746 = ~g744;
  assign g747 = ~g419 | ~g746;
  assign g748 = ~g420 | ~g744;
  assign g749 = ~g747 | ~g748;
  assign g750 = ~g441 & ~g749;
  assign g751 = ~g750;
  assign g752 = ~g441 | ~g749;
  assign g753 = ~g751 | ~g752;
  assign g754 = ~g730 | ~g753;
  assign g755 = ~g753;
  assign g756 = ~g729 | ~g755;
  assign g757 = ~g754 | ~g756;
  assign g758 = ~g757;
  assign g759 = ~g721 | ~g758;
  assign g760 = ~g722 | ~g758;
  assign g761 = ~g721 | ~g757;
  assign g762 = ~g760 | ~g761;
  assign g763 = ~g719 & ~g762;
  assign g764 = ~g719 | ~g762;
  assign g765 = ~g764;
  assign g766 = ~g763 & ~g765;
  assign g767 = ~g759 | ~g764;
  assign g768 = ~g767;
  assign g769 = ~g725 | ~g756;
  assign g770 = ~g745 | ~g752;
  assign g771 = ~g770;
  assign g772 = ~g732 | ~g740;
  assign g773 = ~g736 | ~g772;
  assign g774 = ~g422 | ~g773;
  assign g775 = ~g423 | ~g773;
  assign g776 = ~g773;
  assign g777 = ~g422 | ~g776;
  assign g778 = ~g775 | ~g777;
  assign g779 = ~g778;
  assign g780 = ~g688 | ~g779;
  assign g781 = ~g689 | ~g778;
  assign g782 = ~g780 | ~g781;
  assign g783 = ~g782;
  assign g784 = ~g688 | ~g778;
  assign g785 = ~g774 | ~g784;
  assign g786 = ~g100 | ~g543;
  assign g787 = ~g786;
  assign g788 = ~g348 | ~g787;
  assign g789 = ~g100 | ~g543;
  assign g790 = ~g334 | ~g789;
  assign g791 = ~g788 | ~g790;
  assign g792 = ~g786 | ~g791;
  assign g793 = ~g791;
  assign g794 = ~g787 | ~g793;
  assign g795 = ~g792 | ~g794;
  assign g796 = ~g528 | ~g795;
  assign g797 = ~g795;
  assign g798 = ~g528 | ~g797;
  assign g799 = ~g529 | ~g795;
  assign g800 = ~g798 | ~g799;
  assign g801 = ~g447 & ~g800;
  assign g802 = ~g801;
  assign g803 = ~g447 | ~g800;
  assign g804 = ~g802 | ~g803;
  assign g805 = ~g804;
  assign g806 = ~g782 | ~g805;
  assign g807 = ~g783 | ~g804;
  assign g808 = ~g806 | ~g807;
  assign g809 = ~g770 | ~g808;
  assign g810 = ~g808;
  assign g811 = ~g771 | ~g810;
  assign g812 = ~g809 | ~g811;
  assign g813 = ~g769 & ~g812;
  assign g814 = ~g813;
  assign g815 = ~g769 | ~g812;
  assign g816 = ~g814 | ~g815;
  assign g817 = ~g767 | ~g816;
  assign g818 = ~g816;
  assign g819 = ~g768 | ~g818;
  assign g820 = ~g817 | ~g819;
  assign g821 = ~g767 | ~g818;
  assign g822 = ~g815 | ~g821;
  assign g823 = ~g822;
  assign g824 = ~g770 | ~g810;
  assign g825 = ~g806 | ~g824;
  assign g826 = ~g796 | ~g803;
  assign g827 = ~g826;
  assign g828 = ~g520 | ~g827;
  assign g829 = ~g519 | ~g826;
  assign g830 = ~g828 | ~g829;
  assign g831 = ~g785 & ~g830;
  assign g832 = ~g831;
  assign g833 = ~g785 | ~g830;
  assign g834 = ~g832 | ~g833;
  assign g835 = ~g834;
  assign g836 = ~g520 | ~g826;
  assign g837 = ~g516 | ~g836;
  assign g838 = ~g837;
  assign g839 = ~g786 | ~g793;
  assign g840 = ~g790 | ~g839;
  assign g841 = ~g536 | ~g840;
  assign g842 = ~g840;
  assign g843 = ~g536 | ~g842;
  assign g844 = ~g535 | ~g840;
  assign g845 = ~g843 | ~g844;
  assign g846 = ~g691 & ~g845;
  assign g847 = ~g846;
  assign g848 = ~g691 | ~g845;
  assign g849 = ~g847 | ~g848;
  assign g850 = ~g835 | ~g849;
  assign g851 = ~g849;
  assign g852 = ~g834 | ~g851;
  assign g853 = ~g850 | ~g852;
  assign g854 = ~g825 & ~g853;
  assign g855 = ~g854;
  assign g856 = ~g825 | ~g853;
  assign g857 = ~g855 | ~g856;
  assign g858 = ~g822 | ~g857;
  assign g859 = ~g857;
  assign g860 = ~g823 | ~g859;
  assign g861 = ~g858 | ~g860;
  assign g862 = ~g822 | ~g859;
  assign g863 = ~g856 | ~g862;
  assign g864 = ~g863;
  assign g865 = ~g835 | ~g851;
  assign g866 = ~g833 | ~g865;
  assign g867 = ~g841 | ~g848;
  assign g868 = ~g542 & ~g867;
  assign g869 = ~g868;
  assign g870 = ~g542 | ~g867;
  assign g871 = ~g538 | ~g870;
  assign g872 = ~g507 & ~g871;
  assign g873 = ~g872;
  assign g874 = ~g507 | ~g871;
  assign g875 = ~g505 | ~g874;
  assign g876 = ~g501 & ~g875;
  assign g877 = ~g876;
  assign g878 = ~g501 | ~g875;
  assign g879 = ~g877 | ~g878;
  assign g880 = ~g879;
  assign g881 = ~g873 | ~g874;
  assign g882 = ~g881;
  assign g883 = ~g869 | ~g870;
  assign g884 = ~g883;
  assign g885 = ~g837 | ~g884;
  assign g886 = ~g838 | ~g884;
  assign g887 = ~g837 | ~g883;
  assign g888 = ~g886 | ~g887;
  assign g889 = ~g511 | ~g888;
  assign g890 = ~g885 | ~g889;
  assign g891 = ~g882 | ~g890;
  assign g892 = ~g890;
  assign g893 = ~g882 | ~g892;
  assign g894 = ~g881 | ~g890;
  assign g895 = ~g893 | ~g894;
  assign g896 = ~g888;
  assign g897 = ~g511 | ~g896;
  assign g898 = ~g512 | ~g888;
  assign g899 = ~g897 | ~g898;
  assign g900 = ~g866 & ~g899;
  assign g901 = ~g900;
  assign g902 = ~g866 | ~g899;
  assign g903 = ~g901 | ~g902;
  assign g904 = ~g903;
  assign g905 = ~g863 | ~g904;
  assign g906 = ~g902 | ~g905;
  assign g907 = ~g895 & ~g906;
  assign g908 = ~g895 | ~g906;
  assign g909 = ~g891 | ~g908;
  assign g910 = ~g880 | ~g909;
  assign g911 = ~g878 | ~g910;
  assign g912 = ~g497 & ~g911;
  assign g913 = ~g497 | ~g911;
  assign g914 = ~g493 | ~g913;
  assign g915 = ~g271 | ~g914;
  assign g916 = ~g269 | ~g915;
  assign g917 = ~g215 & ~g916;
  assign g918 = ~g215 | ~g916;
  assign g919 = ~g211 | ~g918;
  assign g920 = 1'b0;
  assign g921 = ~g129 | ~g920;
  assign g922 = ~g921;
  assign g923 = 1'b0;
  assign g924 = ~g133 | ~g923;
  assign g925 = ~g132 | ~g919;
  assign g926 = ~g924 | ~g925;
  assign g927 = ~g918;
  assign g928 = ~g917 & ~g927;
  assign g929 = ~g914;
  assign g930 = ~g271 | ~g929;
  assign g931 = ~g270 | ~g914;
  assign g932 = ~g930 | ~g931;
  assign g933 = ~g913;
  assign g934 = ~g912 & ~g933;
  assign g935 = ~g909;
  assign g936 = ~g880 | ~g935;
  assign g937 = ~g879 | ~g909;
  assign g938 = ~g936 | ~g937;
  assign g939 = ~g908;
  assign g940 = ~g907 & ~g939;
  assign g941 = ~g864 | ~g904;
  assign g942 = ~g863 | ~g903;
  assign g943 = ~g941 | ~g942;
  assign g944 = 1'b0;
  assign g945 = 1'b0;
  assign g946 = g945;
  assign g947 = g550;
  assign g948 = g599;
  assign g949 = g605;
  assign g950 = g634;
  assign g951 = g670;
  assign g952 = g717;
  assign g953 = g766;
  assign g954 = g820;
  assign g955 = g861;
  assign g956 = g943;
  assign g957 = g940;
  assign g958 = g938;
  assign g959 = g934;
  assign g960 = g932;
  assign g961 = g928;
  assign g962 = g926;
  assign g963 = g922;
endmodule


