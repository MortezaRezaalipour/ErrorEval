module adder_i60_o31 (a,b,r);
input [29:0] a,b;
output [30:0] r;

assign r = a+b;

endmodule

