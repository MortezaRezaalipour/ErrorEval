// Benchmark "circuit" written by ABC on Tue Apr 12 01:41:42 2022

module circuit ( 
    g0, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15,
    g16, g17, g18, g19, g20, g21, g22, g23,
    g855, g854, g853, g852, g851, g850, g849, g848, g847, g846, g845, g844,
    g843, g842, g841, g840  );
  input  g0, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14,
    g15, g16, g17, g18, g19, g20, g21, g22, g23;
  output g855, g854, g853, g852, g851, g850, g849, g848, g847, g846, g845,
    g844, g843, g842, g841, g840;
  wire g24, g25, g26, g27, g28, g29, g30, g31, g32, g33, g34, g35, g36, g37,
    g38, g39, g40, g41, g42, g43, g44, g45, g46, g47, g48, g49, g50, g51,
    g52, g53, g54, g55, g56, g57, g58, g59, g60, g61, g62, g63, g64, g65,
    g66, g67, g68, g69, g70, g71, g72, g73, g74, g75, g76, g77, g78, g79,
    g80, g81, g82, g83, g84, g85, g86, g87, g88, g89, g90, g91, g92, g93,
    g94, g95, g96, g97, g98, g99, g100, g101, g102, g103, g104, g105, g106,
    g107, g108, g109, g110, g111, g112, g113, g114, g115, g116, g117, g118,
    g119, g120, g121, g122, g123, g124, g125, g126, g127, g128, g129, g130,
    g131, g132, g133, g134, g135, g136, g137, g138, g139, g140, g141, g142,
    g143, g144, g145, g146, g147, g148, g149, g150, g151, g152, g153, g154,
    g155, g156, g157, g158, g159, g160, g161, g162, g163, g164, g165, g166,
    g167, g168, g169, g170, g171, g172, g173, g174, g175, g176, g177, g178,
    g179, g180, g181, g182, g183, g184, g185, g186, g187, g188, g189, g190,
    g191, g192, g193, g194, g195, g196, g197, g198, g199, g200, g201, g202,
    g203, g204, g205, g206, g207, g208, g209, g210, g211, g212, g213, g214,
    g215, g216, g217, g218, g219, g220, g221, g222, g223, g224, g225, g226,
    g227, g228, g229, g230, g231, g232, g233, g234, g235, g236, g237, g238,
    g239, g240, g241, g242, g243, g244, g245, g246, g247, g248, g249, g250,
    g251, g252, g253, g254, g255, g256, g257, g258, g259, g260, g261, g262,
    g263, g264, g265, g266, g267, g268, g269, g270, g271, g272, g273, g274,
    g275, g276, g277, g278, g279, g280, g281, g282, g283, g284, g285, g286,
    g287, g288, g289, g290, g291, g292, g293, g294, g295, g296, g297, g298,
    g299, g300, g301, g302, g303, g304, g305, g306, g307, g308, g309, g310,
    g311, g312, g313, g314, g315, g316, g317, g318, g319, g320, g321, g322,
    g323, g324, g325, g326, g327, g328, g329, g330, g331, g332, g333, g334,
    g335, g336, g337, g338, g339, g340, g341, g342, g343, g344, g345, g346,
    g347, g348, g349, g350, g351, g352, g353, g354, g355, g356, g357, g358,
    g359, g360, g361, g362, g363, g364, g365, g366, g367, g368, g369, g370,
    g371, g372, g373, g374, g375, g376, g377, g378, g379, g380, g381, g382,
    g383, g384, g385, g386, g387, g388, g389, g390, g391, g392, g393, g394,
    g395, g396, g397, g398, g399, g400, g401, g402, g403, g404, g405, g406,
    g407, g408, g409, g410, g411, g412, g413, g414, g415, g416, g417, g418,
    g419, g420, g421, g422, g423, g424, g425, g426, g427, g428, g429, g430,
    g431, g432, g433, g434, g435, g436, g437, g438, g439, g440, g441, g442,
    g443, g444, g445, g446, g447, g448, g449, g450, g451, g452, g453, g454,
    g455, g456, g457, g458, g459, g460, g461, g462, g463, g464, g465, g466,
    g467, g468, g469, g470, g471, g472, g473, g474, g475, g476, g477, g478,
    g479, g480, g481, g482, g483, g484, g485, g486, g487, g488, g489, g490,
    g491, g492, g493, g494, g495, g496, g497, g498, g499, g500, g501, g502,
    g503, g504, g505, g506, g507, g508, g509, g510, g511, g512, g513, g514,
    g515, g516, g517, g518, g519, g520, g521, g522, g523, g524, g525, g526,
    g527, g528, g529, g530, g531, g532, g533, g534, g535, g536, g537, g538,
    g539, g540, g541, g542, g543, g544, g545, g546, g547, g548, g549, g550,
    g551, g552, g553, g554, g555, g556, g557, g558, g559, g560, g561, g562,
    g563, g564, g565, g566, g567, g568, g569, g570, g571, g572, g573, g574,
    g575, g576, g577, g578, g579, g580, g581, g582, g583, g584, g585, g586,
    g587, g588, g589, g590, g591, g592, g593, g594, g595, g596, g597, g598,
    g599, g600, g601, g602, g603, g604, g605, g606, g607, g608, g609, g610,
    g611, g612, g613, g614, g615, g616, g617, g618, g619, g620, g621, g622,
    g623, g624, g625, g626, g627, g628, g629, g630, g631, g632, g633, g634,
    g635, g636, g637, g638, g639, g640, g641, g642, g643, g644, g645, g646,
    g647, g648, g649, g650, g651, g652, g653, g654, g655, g656, g657, g658,
    g659, g660, g661, g662, g663, g664, g665, g666, g667, g668, g669, g670,
    g671, g672, g673, g674, g675, g676, g677, g678, g679, g680, g681, g682,
    g683, g684, g685, g686, g687, g688, g689, g690, g691, g692, g693, g694,
    g695, g696, g697, g698, g699, g700, g701, g702, g703, g704, g705, g706,
    g707, g708, g709, g710, g711, g712, g713, g714, g715, g716, g717, g718,
    g719, g720, g721, g722, g723, g724, g725, g726, g727, g728, g729, g730,
    g731, g732, g733, g734, g735, g736, g737, g738, g739, g740, g741, g742,
    g743, g744, g745, g746, g747, g748, g749, g750, g751, g752, g753, g754,
    g755, g756, g757, g758, g759, g760, g761, g762, g763, g764, g765, g766,
    g767, g768, g769, g770, g771, g772, g773, g774, g775, g776, g777, g778,
    g779, g780, g781, g782, g783, g784, g785, g786, g787, g788, g789, g790,
    g791, g792, g793, g794, g795, g796, g797, g798, g799, g800, g801, g802,
    g803, g804, g805, g806, g807, g808, g809, g810, g811, g812, g813, g814,
    g815, g816, g817, g818, g819, g820, g821, g822, g823, g824, g825, g826,
    g827, g828, g829, g830, g831, g832, g833, g834, g835, g836;
  assign g24 = 1'b0;
  assign g25 = 1'b0;
  assign g26 = 1'b0;
  assign g27 = 1'b0;
  assign g28 = 1'b0;
  assign g29 = 1'b0;
  assign g30 = 1'b0;
  assign g31 = 1'b0;
  assign g32 = g7 & g15;
  assign g33 = g7 & g14;
  assign g34 = ~g33;
  assign g35 = g7 & g13;
  assign g36 = ~g35;
  assign g37 = g7 & g12;
  assign g38 = g7 & g11;
  assign g39 = ~g38;
  assign g40 = g7 & g10;
  assign g41 = ~g40;
  assign g42 = g7 & g8;
  assign g43 = ~g42;
  assign g44 = g7 & g9;
  assign g45 = ~g44;
  assign g46 = g6 & g15;
  assign g47 = ~g46;
  assign g48 = g33 & g47;
  assign g49 = g33 & g46;
  assign g50 = g34 & g46;
  assign g51 = g48 | g50;
  assign g52 = g6 & g14;
  assign g53 = ~g52;
  assign g54 = g6 & g13;
  assign g55 = ~g54;
  assign g56 = g6 & g12;
  assign g57 = ~g56;
  assign g58 = g38 & g57;
  assign g59 = g38 & g56;
  assign g60 = g39 & g56;
  assign g61 = g58 | g60;
  assign g62 = g6 & g11;
  assign g63 = ~g62;
  assign g64 = g6 & g10;
  assign g65 = ~g64;
  assign g66 = g6 & g8;
  assign g67 = ~g66;
  assign g68 = g6 & g9;
  assign g69 = ~g68;
  assign g70 = g5 & g15;
  assign g71 = ~g70;
  assign g72 = g52 & g71;
  assign g73 = g52 & g70;
  assign g74 = g53 & g70;
  assign g75 = g72 | g74;
  assign g76 = ~g75;
  assign g77 = g35 & g76;
  assign g78 = g35 & g75;
  assign g79 = g73 | g78;
  assign g80 = g51 & g79;
  assign g81 = ~g80;
  assign g82 = g49 | g80;
  assign g83 = g32 & g82;
  assign g84 = ~g83;
  assign g85 = g32 | g82;
  assign g86 = g84 & g85;
  assign g87 = ~g86;
  assign g88 = g51 | g79;
  assign g89 = g81 & g88;
  assign g90 = ~g89;
  assign g91 = g36 & g75;
  assign g92 = g77 | g91;
  assign g93 = g5 & g14;
  assign g94 = ~g93;
  assign g95 = g5 & g13;
  assign g96 = ~g95;
  assign g97 = g5 & g8;
  assign g98 = ~g97;
  assign g99 = g5 & g12;
  assign g100 = ~g99;
  assign g101 = g62 & g100;
  assign g102 = g62 & g99;
  assign g103 = g63 & g99;
  assign g104 = g101 | g103;
  assign g105 = ~g104;
  assign g106 = g40 & g105;
  assign g107 = g40 & g104;
  assign g108 = g102 | g107;
  assign g109 = g41 & g104;
  assign g110 = g106 | g109;
  assign g111 = ~g110;
  assign g112 = g5 & g11;
  assign g113 = ~g112;
  assign g114 = g5 & g9;
  assign g115 = ~g114;
  assign g116 = g5 & g10;
  assign g117 = ~g116;
  assign g118 = g68 & g117;
  assign g119 = g68 & g116;
  assign g120 = ~g119;
  assign g121 = g69 & g116;
  assign g122 = g118 | g121;
  assign g123 = ~g122;
  assign g124 = g4 & g15;
  assign g125 = ~g124;
  assign g126 = g93 & g125;
  assign g127 = g93 & g124;
  assign g128 = g94 & g124;
  assign g129 = g126 | g128;
  assign g130 = ~g129;
  assign g131 = g54 & g130;
  assign g132 = g54 & g129;
  assign g133 = g127 | g132;
  assign g134 = g92 & g133;
  assign g135 = ~g134;
  assign g136 = g92 | g133;
  assign g137 = g135 & g136;
  assign g138 = ~g137;
  assign g139 = g55 & g129;
  assign g140 = g131 | g139;
  assign g141 = g4 & g14;
  assign g142 = ~g141;
  assign g143 = g4 & g8;
  assign g144 = ~g143;
  assign g145 = g4 & g13;
  assign g146 = ~g145;
  assign g147 = g4 & g9;
  assign g148 = ~g147;
  assign g149 = g4 & g11;
  assign g150 = ~g149;
  assign g151 = g4 & g12;
  assign g152 = ~g151;
  assign g153 = g112 & g152;
  assign g154 = g112 & g151;
  assign g155 = g113 & g151;
  assign g156 = g153 | g155;
  assign g157 = ~g156;
  assign g158 = g44 & g157;
  assign g159 = g44 & g156;
  assign g160 = g154 | g159;
  assign g161 = g45 & g156;
  assign g162 = g158 | g161;
  assign g163 = ~g162;
  assign g164 = g4 & g10;
  assign g165 = ~g164;
  assign g166 = g114 & g165;
  assign g167 = g115 & g164;
  assign g168 = g166 | g167;
  assign g169 = g114 & g164;
  assign g170 = ~g169;
  assign g171 = g122 & g170;
  assign g172 = g122 & g169;
  assign g173 = g123 & g169;
  assign g174 = g171 | g173;
  assign g175 = g3 & g15;
  assign g176 = ~g175;
  assign g177 = g141 & g176;
  assign g178 = g141 & g175;
  assign g179 = g142 & g175;
  assign g180 = g177 | g179;
  assign g181 = ~g180;
  assign g182 = g95 & g181;
  assign g183 = g95 & g180;
  assign g184 = g178 | g183;
  assign g185 = g37 & g184;
  assign g186 = ~g185;
  assign g187 = g37 | g184;
  assign g188 = g186 & g187;
  assign g189 = ~g188;
  assign g190 = g96 & g180;
  assign g191 = g182 | g190;
  assign g192 = g108 & g191;
  assign g193 = ~g192;
  assign g194 = g108 | g191;
  assign g195 = g193 & g194;
  assign g196 = ~g195;
  assign g197 = g3 & g8;
  assign g198 = ~g197;
  assign g199 = g3 & g9;
  assign g200 = ~g199;
  assign g201 = g3 & g14;
  assign g202 = ~g201;
  assign g203 = g3 & g12;
  assign g204 = ~g203;
  assign g205 = g42 & g204;
  assign g206 = g42 & g203;
  assign g207 = g43 & g203;
  assign g208 = g205 | g207;
  assign g209 = ~g208;
  assign g210 = g3 & g11;
  assign g211 = ~g210;
  assign g212 = g3 & g10;
  assign g213 = ~g212;
  assign g214 = g147 & g213;
  assign g215 = g148 & g212;
  assign g216 = g214 | g215;
  assign g217 = ~g216;
  assign g218 = g147 & g212;
  assign g219 = ~g218;
  assign g220 = g3 & g13;
  assign g221 = ~g220;
  assign g222 = g2 & g8;
  assign g223 = ~g222;
  assign g224 = g2 & g9;
  assign g225 = ~g224;
  assign g226 = g2 & g10;
  assign g227 = ~g226;
  assign g228 = g199 & g227;
  assign g229 = g200 & g226;
  assign g230 = g228 | g229;
  assign g231 = ~g230;
  assign g232 = g199 & g226;
  assign g233 = ~g232;
  assign g234 = g97 & g233;
  assign g235 = g97 & g232;
  assign g236 = g98 & g232;
  assign g237 = g234 | g236;
  assign g238 = ~g237;
  assign g239 = g216 & g238;
  assign g240 = g217 & g237;
  assign g241 = g239 | g240;
  assign g242 = ~g241;
  assign g243 = g216 & g237;
  assign g244 = g235 | g243;
  assign g245 = ~g244;
  assign g246 = g2 & g11;
  assign g247 = ~g246;
  assign g248 = g2 & g15;
  assign g249 = ~g248;
  assign g250 = g201 & g249;
  assign g251 = g201 & g248;
  assign g252 = g202 & g248;
  assign g253 = g250 | g252;
  assign g254 = ~g253;
  assign g255 = g145 & g254;
  assign g256 = g145 & g253;
  assign g257 = g251 | g256;
  assign g258 = g61 & g257;
  assign g259 = ~g258;
  assign g260 = g59 | g258;
  assign g261 = ~g260;
  assign g262 = g188 & g261;
  assign g263 = g188 & g260;
  assign g264 = g185 | g263;
  assign g265 = ~g264;
  assign g266 = g137 & g265;
  assign g267 = g137 & g264;
  assign g268 = g134 | g267;
  assign g269 = ~g268;
  assign g270 = g89 & g269;
  assign g271 = g89 & g268;
  assign g272 = g90 & g268;
  assign g273 = g270 | g272;
  assign g274 = g138 & g264;
  assign g275 = g266 | g274;
  assign g276 = g189 & g260;
  assign g277 = g262 | g276;
  assign g278 = g61 | g257;
  assign g279 = g259 & g278;
  assign g280 = ~g279;
  assign g281 = g146 & g253;
  assign g282 = g255 | g281;
  assign g283 = ~g282;
  assign g284 = g110 & g283;
  assign g285 = g110 & g282;
  assign g286 = g111 & g282;
  assign g287 = g284 | g286;
  assign g288 = g2 & g13;
  assign g289 = ~g288;
  assign g290 = g208 & g289;
  assign g291 = g208 & g288;
  assign g292 = g206 | g291;
  assign g293 = ~g292;
  assign g294 = g209 & g288;
  assign g295 = g290 | g294;
  assign g296 = g2 & g12;
  assign g297 = ~g296;
  assign g298 = g210 & g297;
  assign g299 = g210 & g296;
  assign g300 = g211 & g296;
  assign g301 = g298 | g300;
  assign g302 = ~g301;
  assign g303 = g218 & g302;
  assign g304 = g219 & g301;
  assign g305 = g303 | g304;
  assign g306 = ~g305;
  assign g307 = g218 & g301;
  assign g308 = g299 | g307;
  assign g309 = g295 & g308;
  assign g310 = ~g309;
  assign g311 = g295 | g308;
  assign g312 = g310 & g311;
  assign g313 = g2 & g14;
  assign g314 = ~g313;
  assign g315 = g220 & g314;
  assign g316 = g220 & g313;
  assign g317 = g221 & g313;
  assign g318 = g315 | g317;
  assign g319 = ~g318;
  assign g320 = g119 & g319;
  assign g321 = g119 & g318;
  assign g322 = g316 | g321;
  assign g323 = ~g322;
  assign g324 = g120 & g318;
  assign g325 = g320 | g324;
  assign g326 = ~g325;
  assign g327 = g162 & g326;
  assign g328 = g162 & g325;
  assign g329 = g163 & g325;
  assign g330 = g327 | g329;
  assign g331 = g1 & g8;
  assign g332 = ~g331;
  assign g333 = g1 & g9;
  assign g334 = ~g333;
  assign g335 = g1 & g10;
  assign g336 = ~g335;
  assign g337 = g198 | g336;
  assign g338 = g1 & g11;
  assign g339 = ~g338;
  assign g340 = g1 & g12;
  assign g341 = ~g340;
  assign g342 = g1 & g15;
  assign g343 = ~g342;
  assign g344 = g64 & g343;
  assign g345 = g64 & g342;
  assign g346 = g160 | g345;
  assign g347 = g160 & g345;
  assign g348 = ~g347;
  assign g349 = g346 & g348;
  assign g350 = ~g349;
  assign g351 = g322 & g350;
  assign g352 = g322 & g349;
  assign g353 = g323 & g349;
  assign g354 = g351 | g353;
  assign g355 = g347 | g352;
  assign g356 = ~g355;
  assign g357 = g195 & g356;
  assign g358 = g195 & g355;
  assign g359 = g192 | g358;
  assign g360 = g140 & g359;
  assign g361 = ~g360;
  assign g362 = g140 | g359;
  assign g363 = g361 & g362;
  assign g364 = g277 & g363;
  assign g365 = ~g364;
  assign g366 = g360 | g364;
  assign g367 = g275 & g366;
  assign g368 = ~g367;
  assign g369 = g275 | g366;
  assign g370 = g368 & g369;
  assign g371 = ~g370;
  assign g372 = g277 | g363;
  assign g373 = g365 & g372;
  assign g374 = ~g373;
  assign g375 = g196 & g355;
  assign g376 = g357 | g375;
  assign g377 = ~g376;
  assign g378 = g65 & g342;
  assign g379 = g344 | g378;
  assign g380 = g1 & g14;
  assign g381 = ~g380;
  assign g382 = g1 & g13;
  assign g383 = ~g382;
  assign g384 = g0 & g9;
  assign g385 = ~g384;
  assign g386 = g331 & g385;
  assign g387 = g332 & g384;
  assign g388 = g386 | g387;
  assign g389 = 1'b0;
  assign g390 = 1'b0;
  assign g391 = 1'b0;
  assign g392 = 1'b0;
  assign g393 = 1'b0;
  assign g394 = g331 & g384;
  assign g395 = ~g394;
  assign g396 = g0 & g10;
  assign g397 = ~g396;
  assign g398 = g333 & g397;
  assign g399 = g334 & g396;
  assign g400 = g398 | g399;
  assign g401 = ~g400;
  assign g402 = g222 & g401;
  assign g403 = g222 & g400;
  assign g404 = g223 & g400;
  assign g405 = g402 | g404;
  assign g406 = ~g405;
  assign g407 = g394 & g406;
  assign g408 = g395 & g405;
  assign g409 = g407 | g408;
  assign g410 = 1'b0;
  assign g411 = 1'b0;
  assign g412 = 1'b0;
  assign g413 = 1'b0;
  assign g414 = g394 & g405;
  assign g415 = g403 | g414;
  assign g416 = g333 & g396;
  assign g417 = ~g416;
  assign g418 = g197 & g417;
  assign g419 = g337 & g417;
  assign g420 = ~g419;
  assign g421 = g198 & g416;
  assign g422 = g418 | g421;
  assign g423 = ~g422;
  assign g424 = g335 & g423;
  assign g425 = g336 & g422;
  assign g426 = g424 | g425;
  assign g427 = ~g426;
  assign g428 = g0 & g11;
  assign g429 = ~g428;
  assign g430 = g224 & g429;
  assign g431 = g225 & g428;
  assign g432 = g430 | g431;
  assign g433 = ~g432;
  assign g434 = g426 & g433;
  assign g435 = g426 & g432;
  assign g436 = g427 & g432;
  assign g437 = g434 | g436;
  assign g438 = g415 | g437;
  assign g439 = g415 & g437;
  assign g440 = ~g439;
  assign g441 = g438 & g440;
  assign g442 = 1'b0;
  assign g443 = 1'b0;
  assign g444 = 1'b0;
  assign g445 = 1'b0;
  assign g446 = g435 | g439;
  assign g447 = ~g446;
  assign g448 = g224 & g428;
  assign g449 = ~g448;
  assign g450 = g230 & g449;
  assign g451 = g230 & g448;
  assign g452 = g231 & g448;
  assign g453 = g450 | g452;
  assign g454 = ~g453;
  assign g455 = g419 & g454;
  assign g456 = g420 & g453;
  assign g457 = g455 | g456;
  assign g458 = ~g457;
  assign g459 = g451 | g456;
  assign g460 = ~g459;
  assign g461 = g0 & g12;
  assign g462 = ~g461;
  assign g463 = g338 & g462;
  assign g464 = g338 & g461;
  assign g465 = g339 & g461;
  assign g466 = g463 | g465;
  assign g467 = ~g466;
  assign g468 = g143 & g467;
  assign g469 = g144 & g466;
  assign g470 = g468 | g469;
  assign g471 = ~g470;
  assign g472 = g457 & g471;
  assign g473 = g458 & g470;
  assign g474 = g472 | g473;
  assign g475 = ~g474;
  assign g476 = g447 & g475;
  assign g477 = g446 & g475;
  assign g478 = g473 | g477;
  assign g479 = g446 & g474;
  assign g480 = g476 | g479;
  assign g481 = 1'b0;
  assign g482 = 1'b0;
  assign g483 = 1'b0;
  assign g484 = 1'b0;
  assign g485 = g143 & g466;
  assign g486 = g464 | g485;
  assign g487 = g0 & g13;
  assign g488 = ~g487;
  assign g489 = g340 & g488;
  assign g490 = g340 & g487;
  assign g491 = g341 & g487;
  assign g492 = g489 | g491;
  assign g493 = ~g492;
  assign g494 = g246 & g493;
  assign g495 = g247 & g492;
  assign g496 = g494 | g495;
  assign g497 = g486 & g496;
  assign g498 = ~g497;
  assign g499 = g486 | g496;
  assign g500 = g498 & g499;
  assign g501 = ~g500;
  assign g502 = g459 & g501;
  assign g503 = g460 & g500;
  assign g504 = g502 | g503;
  assign g505 = ~g504;
  assign g506 = g241 & g505;
  assign g507 = g241 & g504;
  assign g508 = g242 & g504;
  assign g509 = g506 | g508;
  assign g510 = g478 | g509;
  assign g511 = g478 & g509;
  assign g512 = ~g511;
  assign g513 = g510 & g512;
  assign g514 = 1'b0;
  assign g515 = 1'b0;
  assign g516 = 1'b0;
  assign g517 = 1'b0;
  assign g518 = g507 | g511;
  assign g519 = ~g518;
  assign g520 = g459 & g500;
  assign g521 = g497 | g520;
  assign g522 = g246 & g492;
  assign g523 = g490 | g522;
  assign g524 = g168 & g523;
  assign g525 = ~g524;
  assign g526 = g168 | g523;
  assign g527 = g525 & g526;
  assign g528 = ~g527;
  assign g529 = g244 & g528;
  assign g530 = g245 & g527;
  assign g531 = g529 | g530;
  assign g532 = g244 & g527;
  assign g533 = g524 | g532;
  assign g534 = ~g533;
  assign g535 = g0 & g15;
  assign g536 = ~g535;
  assign g537 = g380 & g536;
  assign g538 = g380 & g535;
  assign g539 = g381 & g535;
  assign g540 = g537 | g539;
  assign g541 = ~g540;
  assign g542 = g149 & g541;
  assign g543 = g149 & g540;
  assign g544 = g538 | g543;
  assign g545 = g379 & g544;
  assign g546 = ~g545;
  assign g547 = g379 | g544;
  assign g548 = g546 & g547;
  assign g549 = ~g548;
  assign g550 = g292 & g549;
  assign g551 = g292 & g548;
  assign g552 = g545 | g551;
  assign g553 = g287 & g552;
  assign g554 = ~g553;
  assign g555 = g285 | g553;
  assign g556 = ~g555;
  assign g557 = g279 & g556;
  assign g558 = g279 & g555;
  assign g559 = g280 & g555;
  assign g560 = g557 | g559;
  assign g561 = ~g560;
  assign g562 = g376 & g561;
  assign g563 = g376 & g560;
  assign g564 = g558 | g563;
  assign g565 = ~g564;
  assign g566 = g373 & g565;
  assign g567 = g373 & g564;
  assign g568 = g374 & g564;
  assign g569 = g566 | g568;
  assign g570 = g377 & g560;
  assign g571 = g562 | g570;
  assign g572 = g287 | g552;
  assign g573 = g554 & g572;
  assign g574 = ~g573;
  assign g575 = g293 & g548;
  assign g576 = g550 | g575;
  assign g577 = g150 & g540;
  assign g578 = g542 | g577;
  assign g579 = g312 | g578;
  assign g580 = g312 & g578;
  assign g581 = ~g580;
  assign g582 = g579 & g581;
  assign g583 = ~g582;
  assign g584 = g309 | g580;
  assign g585 = g576 & g584;
  assign g586 = ~g585;
  assign g587 = g576 | g584;
  assign g588 = g586 & g587;
  assign g589 = ~g588;
  assign g590 = g0 & g14;
  assign g591 = ~g590;
  assign g592 = g382 & g591;
  assign g593 = g382 & g590;
  assign g594 = g383 & g590;
  assign g595 = g592 | g594;
  assign g596 = ~g595;
  assign g597 = g66 & g596;
  assign g598 = g67 & g595;
  assign g599 = g597 | g598;
  assign g600 = ~g599;
  assign g601 = g305 & g600;
  assign g602 = g305 & g599;
  assign g603 = g306 & g599;
  assign g604 = g601 | g603;
  assign g605 = g521 | g604;
  assign g606 = g521 & g604;
  assign g607 = ~g606;
  assign g608 = g605 & g607;
  assign g609 = g531 & g608;
  assign g610 = ~g609;
  assign g611 = g531 | g608;
  assign g612 = g610 & g611;
  assign g613 = ~g612;
  assign g614 = g518 & g613;
  assign g615 = g519 & g612;
  assign g616 = g614 | g615;
  assign g617 = 1'b0;
  assign g618 = 1'b0;
  assign g619 = 1'b0;
  assign g620 = 1'b0;
  assign g621 = g518 & g612;
  assign g622 = g609 | g621;
  assign g623 = g602 | g606;
  assign g624 = g66 & g595;
  assign g625 = g593 | g624;
  assign g626 = g174 | g625;
  assign g627 = g174 & g625;
  assign g628 = ~g627;
  assign g629 = g626 & g628;
  assign g630 = ~g629;
  assign g631 = g533 & g630;
  assign g632 = g533 & g629;
  assign g633 = g534 & g629;
  assign g634 = g631 | g633;
  assign g635 = g623 | g634;
  assign g636 = g623 & g634;
  assign g637 = ~g636;
  assign g638 = g635 & g637;
  assign g639 = ~g638;
  assign g640 = g582 & g639;
  assign g641 = g582 & g638;
  assign g642 = g583 & g638;
  assign g643 = g640 | g642;
  assign g644 = g622 | g643;
  assign g645 = g622 & g643;
  assign g646 = ~g645;
  assign g647 = g644 & g646;
  assign g648 = 1'b0;
  assign g649 = 1'b0;
  assign g650 = 1'b0;
  assign g651 = 1'b0;
  assign g652 = g641 | g645;
  assign g653 = ~g652;
  assign g654 = g632 | g636;
  assign g655 = g172 | g627;
  assign g656 = g330 & g655;
  assign g657 = ~g656;
  assign g658 = g328 | g656;
  assign g659 = g354 & g658;
  assign g660 = ~g659;
  assign g661 = g354 | g658;
  assign g662 = g660 & g661;
  assign g663 = ~g662;
  assign g664 = g573 & g663;
  assign g665 = g573 & g662;
  assign g666 = g659 | g665;
  assign g667 = g571 & g666;
  assign g668 = ~g667;
  assign g669 = g571 | g666;
  assign g670 = g668 & g669;
  assign g671 = ~g670;
  assign g672 = g574 & g662;
  assign g673 = g664 | g672;
  assign g674 = g330 | g655;
  assign g675 = g657 & g674;
  assign g676 = ~g675;
  assign g677 = g588 & g676;
  assign g678 = g589 & g675;
  assign g679 = g677 | g678;
  assign g680 = g654 & g679;
  assign g681 = ~g680;
  assign g682 = g654 | g679;
  assign g683 = g681 & g682;
  assign g684 = ~g683;
  assign g685 = g652 & g684;
  assign g686 = g653 & g683;
  assign g687 = g685 | g686;
  assign g688 = g652 & g683;
  assign g689 = g680 | g688;
  assign g690 = ~g689;
  assign g691 = g588 & g675;
  assign g692 = g585 | g691;
  assign g693 = g673 & g692;
  assign g694 = ~g693;
  assign g695 = g673 | g692;
  assign g696 = g694 & g695;
  assign g697 = ~g696;
  assign g698 = g689 & g697;
  assign g699 = g690 & g696;
  assign g700 = g698 | g699;
  assign g701 = 1'b0;
  assign g702 = g689 & g696;
  assign g703 = g693 | g702;
  assign g704 = ~g703;
  assign g705 = g670 & g704;
  assign g706 = g670 & g703;
  assign g707 = g667 | g706;
  assign g708 = g569 | g707;
  assign g709 = g569 & g707;
  assign g710 = ~g709;
  assign g711 = g708 & g710;
  assign g712 = 1'b0;
  assign g713 = g567 | g709;
  assign g714 = ~g713;
  assign g715 = g370 & g714;
  assign g716 = g370 & g713;
  assign g717 = g367 | g716;
  assign g718 = g273 | g717;
  assign g719 = g273 & g717;
  assign g720 = ~g719;
  assign g721 = g718 & g720;
  assign g722 = 1'b0;
  assign g723 = g271 | g719;
  assign g724 = ~g723;
  assign g725 = g86 & g724;
  assign g726 = g86 & g723;
  assign g727 = g83 | g726;
  assign g728 = ~g727;
  assign g729 = g87 & g723;
  assign g730 = g725 | g729;
  assign g731 = 1'b0;
  assign g732 = g371 & g713;
  assign g733 = g715 | g732;
  assign g734 = 1'b0;
  assign g735 = g671 & g703;
  assign g736 = g705 | g735;
  assign g737 = 1'b0;
  assign g738 = g0 & g8;
  assign g739 = 1'b0;
  assign g740 = 1'b0;
  assign g741 = g16 & g738;
  assign g742 = 1'b0;
  assign g743 = 1'b0;
  assign g744 = 1'b0;
  assign g745 = 1'b0;
  assign g746 = g388 & g741;
  assign g747 = g388 | g741;
  assign g748 = g17 & g747;
  assign g749 = g746 | g748;
  assign g750 = 1'b0;
  assign g751 = 1'b0;
  assign g752 = 1'b0;
  assign g753 = 1'b0;
  assign g754 = g409 & g749;
  assign g755 = g409 | g749;
  assign g756 = g18 & g755;
  assign g757 = g754 | g756;
  assign g758 = 1'b0;
  assign g759 = 1'b0;
  assign g760 = 1'b0;
  assign g761 = 1'b0;
  assign g762 = g441 & g757;
  assign g763 = g441 | g757;
  assign g764 = g19 & g763;
  assign g765 = g762 | g764;
  assign g766 = 1'b0;
  assign g767 = 1'b0;
  assign g768 = 1'b0;
  assign g769 = 1'b0;
  assign g770 = g480 & g765;
  assign g771 = g480 | g765;
  assign g772 = g20 & g771;
  assign g773 = g770 | g772;
  assign g774 = 1'b0;
  assign g775 = 1'b0;
  assign g776 = 1'b0;
  assign g777 = 1'b0;
  assign g778 = g513 & g773;
  assign g779 = g513 | g773;
  assign g780 = g21 & g779;
  assign g781 = g778 | g780;
  assign g782 = 1'b0;
  assign g783 = 1'b0;
  assign g784 = 1'b0;
  assign g785 = 1'b0;
  assign g786 = g616 & g781;
  assign g787 = g616 | g781;
  assign g788 = g22 & g787;
  assign g789 = g786 | g788;
  assign g790 = 1'b0;
  assign g791 = 1'b0;
  assign g792 = 1'b0;
  assign g793 = 1'b0;
  assign g794 = g647 & g789;
  assign g795 = g647 | g789;
  assign g796 = g23 & g795;
  assign g797 = g794 | g796;
  assign g798 = 1'b0;
  assign g799 = g687 & g797;
  assign g800 = 1'b0;
  assign g801 = 1'b0;
  assign g802 = 1'b0;
  assign g803 = 1'b0;
  assign g804 = 1'b0;
  assign g805 = g700 & g799;
  assign g806 = 1'b0;
  assign g807 = 1'b0;
  assign g808 = g736 & g805;
  assign g809 = 1'b0;
  assign g810 = 1'b0;
  assign g811 = g711 & g808;
  assign g812 = 1'b0;
  assign g813 = 1'b0;
  assign g814 = g733 & g811;
  assign g815 = 1'b0;
  assign g816 = 1'b0;
  assign g817 = g721 & g814;
  assign g818 = 1'b0;
  assign g819 = 1'b0;
  assign g820 = g730 & g817;
  assign g821 = ~g820;
  assign g822 = g727 & g821;
  assign g823 = g728 & g820;
  assign g824 = g822 | g823;
  assign g825 = 1'b0;
  assign g826 = 1'b0;
  assign g827 = 1'b0;
  assign g828 = 1'b0;
  assign g829 = 1'b0;
  assign g830 = 1'b0;
  assign g831 = 1'b0;
  assign g832 = 1'b0;
  assign g833 = 1'b0;
  assign g834 = 1'b0;
  assign g835 = 1'b0;
  assign g836 = 1'b0;
  assign g840 = g836;
  assign g841 = g745;
  assign g842 = g753;
  assign g843 = g761;
  assign g844 = g769;
  assign g845 = g777;
  assign g846 = g785;
  assign g847 = g793;
  assign g848 = g802;
  assign g849 = g804;
  assign g850 = g834;
  assign g851 = g832;
  assign g852 = g830;
  assign g853 = g828;
  assign g854 = g826;
  assign g855 = g824;
endmodule


