module top(pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, po0, po1, po2, po3, po4, po5);
  input pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8;
  output po0, po1, po2, po3, po4, po5;
  wire n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70;
  assign n10 = pi0 & pi3;
  assign n11 = pi6 & n10;
  assign n12 = ~pi6 & ~n10;
  assign n13 = ~n11 & ~n12;
  assign n14 = pi0 & pi4;
  assign n15 = pi1 & pi3;
  assign n16 = pi7 & n15;
  assign n17 = ~pi7 & ~n15;
  assign n18 = ~n16 & ~n17;
  assign n19 = n14 & n18;
  assign n20 = ~n14 & ~n18;
  assign n21 = ~n19 & ~n20;
  assign n22 = n11 & n21;
  assign n23 = ~n11 & ~n21;
  assign n24 = ~n22 & ~n23;
  assign n25 = pi0 & pi5;
  assign n26 = ~n16 & ~n19;
  assign n27 = pi1 & pi4;
  assign n28 = pi2 & pi3;
  assign n29 = pi8 & n28;
  assign n30 = ~pi8 & ~n28;
  assign n31 = ~n29 & ~n30;
  assign n32 = n27 & n31;
  assign n33 = ~n27 & ~n31;
  assign n34 = ~n32 & ~n33;
  assign n35 = ~n26 & n34;
  assign n36 = n26 & ~n34;
  assign n37 = ~n35 & ~n36;
  assign n38 = n25 & n37;
  assign n39 = ~n25 & ~n37;
  assign n40 = ~n38 & ~n39;
  assign n41 = n22 & n40;
  assign n42 = ~n22 & ~n40;
  assign n43 = ~n41 & ~n42;
  assign n44 = ~n35 & ~n38;
  assign n45 = ~n29 & ~n32;
  assign n46 = pi2 & pi5;
  assign n47 = n27 & n46;
  assign n48 = pi1 & pi5;
  assign n49 = pi2 & pi4;
  assign n50 = ~n48 & ~n49;
  assign n51 = ~n47 & ~n50;
  assign n52 = ~n45 & n51;
  assign n53 = n45 & ~n51;
  assign n54 = ~n52 & ~n53;
  assign n55 = ~n44 & n54;
  assign n56 = n44 & ~n54;
  assign n57 = ~n55 & ~n56;
  assign n58 = n41 & n57;
  assign n59 = ~n41 & ~n57;
  assign n60 = ~n58 & ~n59;
  assign n61 = ~n55 & ~n58;
  assign n62 = ~n27 & n46;
  assign n63 = n52 & n62;
  assign n64 = ~n52 & ~n62;
  assign n65 = ~n63 & ~n64;
  assign n66 = ~n61 & n65;
  assign n67 = n61 & ~n65;
  assign n68 = ~n66 & ~n67;
  assign n69 = ~n47 & ~n63;
  assign n70 = ~n66 & n69;
  assign po0 = n13;
  assign po1 = n24;
  assign po2 = n43;
  assign po3 = n60;
  assign po4 = n68;
  assign po5 = ~n70;
endmodule
