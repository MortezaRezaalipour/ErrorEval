module madd_8_app3(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15;
  wire n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536;
  assign n25 = pi00 & pi09;
  assign n26 = pi02 & pi11;
  assign n27 = n25 & n26;
  assign n28 = pi00 & pi11;
  assign n29 = pi02 & pi09;
  assign n30 = ~n28 & ~n29;
  assign n31 = ~n27 & ~n30;
  assign n32 = pi03 & pi08;
  assign n33 = pi01 & pi10;
  assign n34 = ~n25 & n33;
  assign n35 = n32 & ~n34;
  assign n36 = ~n32 & n34;
  assign n37 = ~n35 & ~n36;
  assign n38 = n31 & ~n37;
  assign n39 = ~n31 & n37;
  assign n40 = ~n38 & ~n39;
  assign n41 = pi02 & pi08;
  assign n42 = pi00 & pi10;
  assign n43 = pi01 & pi09;
  assign n44 = n42 & ~n43;
  assign n45 = ~n42 & n43;
  assign n46 = ~n44 & ~n45;
  assign n47 = n41 & ~n46;
  assign n48 = pi00 & pi08;
  assign n49 = n43 & n48;
  assign n50 = ~n42 & ~n43;
  assign n51 = n25 & n33;
  assign n52 = ~n50 & ~n51;
  assign n53 = ~n41 & ~n52;
  assign n54 = ~n47 & ~n53;
  assign n55 = n49 & n54;
  assign n56 = ~n47 & ~n55;
  assign n57 = ~n40 & n56;
  assign n58 = n40 & ~n56;
  assign n59 = ~n57 & ~n58;
  assign n60 = pi16 & n48;
  assign n61 = ~pi17 & ~n60;
  assign n62 = pi17 & n60;
  assign n63 = pi01 & pi08;
  assign n64 = ~n25 & ~n63;
  assign n65 = ~n49 & ~n64;
  assign n66 = ~n62 & ~n65;
  assign n67 = ~n61 & ~n66;
  assign n68 = ~pi18 & ~n67;
  assign n69 = ~n61 & n65;
  assign n70 = ~n62 & ~n69;
  assign n71 = pi18 & ~n70;
  assign n72 = ~n49 & ~n54;
  assign n73 = ~n55 & ~n72;
  assign n74 = ~n71 & ~n73;
  assign n75 = ~n68 & ~n74;
  assign n76 = ~n59 & ~n75;
  assign n77 = ~n68 & n73;
  assign n78 = ~n71 & ~n77;
  assign n79 = n59 & ~n78;
  assign n80 = ~pi19 & ~n79;
  assign n81 = ~n76 & ~n80;
  assign n82 = pi01 & pi12;
  assign n83 = n28 & n82;
  assign n84 = pi00 & pi12;
  assign n85 = pi01 & pi11;
  assign n86 = ~n84 & ~n85;
  assign n87 = ~n83 & ~n86;
  assign n88 = pi04 & pi08;
  assign n89 = n87 & n88;
  assign n90 = ~n87 & ~n88;
  assign n91 = ~n89 & ~n90;
  assign n92 = pi03 & pi10;
  assign n93 = n29 & n92;
  assign n94 = pi02 & pi10;
  assign n95 = pi03 & pi09;
  assign n96 = ~n94 & ~n95;
  assign n97 = ~n93 & ~n96;
  assign n98 = n27 & n97;
  assign n99 = ~n27 & ~n97;
  assign n100 = ~n98 & ~n99;
  assign n101 = ~n25 & ~n32;
  assign n102 = n33 & ~n101;
  assign n103 = n100 & n102;
  assign n104 = ~n100 & ~n102;
  assign n105 = ~n103 & ~n104;
  assign n106 = n91 & n105;
  assign n107 = ~n91 & ~n105;
  assign n108 = ~n106 & ~n107;
  assign n109 = ~n38 & ~n58;
  assign n110 = n108 & ~n109;
  assign n111 = ~n108 & n109;
  assign n112 = ~n110 & ~n111;
  assign n113 = ~n81 & ~n112;
  assign n114 = pi19 & ~n76;
  assign n115 = ~n79 & ~n114;
  assign n116 = n112 & ~n115;
  assign n117 = ~pi20 & ~n116;
  assign n118 = ~n113 & ~n117;
  assign n119 = pi00 & pi13;
  assign n120 = ~n82 & ~n119;
  assign n121 = n82 & n119;
  assign n122 = ~n120 & ~n121;
  assign n123 = n26 & n122;
  assign n124 = ~n26 & ~n122;
  assign n125 = ~n123 & ~n124;
  assign n126 = ~n83 & ~n89;
  assign n127 = ~n125 & n126;
  assign n128 = n125 & ~n126;
  assign n129 = ~n127 & ~n128;
  assign n130 = ~n98 & ~n103;
  assign n131 = n129 & ~n130;
  assign n132 = ~n129 & n130;
  assign n133 = ~n131 & ~n132;
  assign n134 = pi05 & pi08;
  assign n135 = n93 & n134;
  assign n136 = ~n93 & ~n134;
  assign n137 = ~n135 & ~n136;
  assign n138 = pi04 & pi09;
  assign n139 = n92 & n138;
  assign n140 = ~n92 & ~n138;
  assign n141 = ~n139 & ~n140;
  assign n142 = n137 & n141;
  assign n143 = ~n137 & ~n141;
  assign n144 = ~n142 & ~n143;
  assign n145 = n133 & n144;
  assign n146 = ~n133 & ~n144;
  assign n147 = ~n145 & ~n146;
  assign n148 = ~n106 & ~n110;
  assign n149 = n147 & ~n148;
  assign n150 = ~n147 & n148;
  assign n151 = ~n149 & ~n150;
  assign n152 = ~n118 & ~n151;
  assign n153 = pi20 & ~n113;
  assign n154 = ~n116 & ~n153;
  assign n155 = n151 & ~n154;
  assign n156 = ~pi21 & ~n155;
  assign n157 = ~n152 & ~n156;
  assign n158 = ~n135 & ~n142;
  assign n159 = ~n121 & ~n123;
  assign n160 = pi05 & pi10;
  assign n161 = n138 & n160;
  assign n162 = pi04 & pi10;
  assign n163 = pi05 & pi09;
  assign n164 = ~n162 & ~n163;
  assign n165 = ~n161 & ~n164;
  assign n166 = ~n159 & n165;
  assign n167 = n159 & ~n165;
  assign n168 = ~n166 & ~n167;
  assign n169 = ~n158 & n168;
  assign n170 = n158 & ~n168;
  assign n171 = ~n169 & ~n170;
  assign n172 = pi01 & pi13;
  assign n173 = pi00 & pi14;
  assign n174 = ~n172 & ~n173;
  assign n175 = pi01 & pi14;
  assign n176 = n119 & n175;
  assign n177 = ~n174 & ~n176;
  assign n178 = pi06 & pi08;
  assign n179 = n177 & n178;
  assign n180 = ~n177 & ~n178;
  assign n181 = ~n179 & ~n180;
  assign n182 = pi02 & pi12;
  assign n183 = pi03 & pi11;
  assign n184 = ~n182 & ~n183;
  assign n185 = pi03 & pi12;
  assign n186 = n26 & n185;
  assign n187 = ~n184 & ~n186;
  assign n188 = n139 & n187;
  assign n189 = ~n139 & ~n187;
  assign n190 = ~n188 & ~n189;
  assign n191 = n181 & n190;
  assign n192 = ~n181 & ~n190;
  assign n193 = ~n191 & ~n192;
  assign n194 = ~n128 & ~n131;
  assign n195 = n193 & ~n194;
  assign n196 = ~n193 & n194;
  assign n197 = ~n195 & ~n196;
  assign n198 = ~n171 & ~n197;
  assign n199 = n171 & n197;
  assign n200 = ~n198 & ~n199;
  assign n201 = ~n145 & ~n149;
  assign n202 = n200 & ~n201;
  assign n203 = ~n200 & n201;
  assign n204 = ~n202 & ~n203;
  assign n205 = ~n157 & ~n204;
  assign n206 = pi21 & ~n152;
  assign n207 = ~n155 & ~n206;
  assign n208 = n204 & ~n207;
  assign n209 = ~pi22 & ~n208;
  assign n210 = ~n205 & ~n209;
  assign n211 = ~n166 & ~n169;
  assign n212 = ~n176 & ~n179;
  assign n213 = pi06 & pi09;
  assign n214 = ~n138 & n160;
  assign n215 = n213 & ~n214;
  assign n216 = ~n213 & n214;
  assign n217 = ~n215 & ~n216;
  assign n218 = ~n212 & ~n217;
  assign n219 = ~n213 & ~n214;
  assign n220 = n213 & n214;
  assign n221 = ~n219 & ~n220;
  assign n222 = n212 & ~n221;
  assign n223 = ~n218 & ~n222;
  assign n224 = n211 & ~n223;
  assign n225 = ~n211 & n223;
  assign n226 = ~n224 & ~n225;
  assign n227 = ~n191 & ~n195;
  assign n228 = ~n226 & n227;
  assign n229 = n226 & ~n227;
  assign n230 = ~n228 & ~n229;
  assign n231 = pi00 & pi15;
  assign n232 = ~n175 & ~n231;
  assign n233 = n175 & n231;
  assign n234 = ~n232 & ~n233;
  assign n235 = pi04 & pi11;
  assign n236 = n234 & n235;
  assign n237 = ~n234 & ~n235;
  assign n238 = ~n236 & ~n237;
  assign n239 = ~n186 & ~n188;
  assign n240 = pi02 & pi13;
  assign n241 = pi07 & pi12;
  assign n242 = n32 & n241;
  assign n243 = pi07 & pi08;
  assign n244 = ~n185 & ~n243;
  assign n245 = ~n242 & ~n244;
  assign n246 = ~n240 & ~n245;
  assign n247 = n240 & n245;
  assign n248 = ~n246 & ~n247;
  assign n249 = ~n239 & n248;
  assign n250 = n239 & ~n248;
  assign n251 = ~n249 & ~n250;
  assign n252 = n238 & n251;
  assign n253 = ~n238 & ~n251;
  assign n254 = ~n252 & ~n253;
  assign n255 = n230 & n254;
  assign n256 = ~n230 & ~n254;
  assign n257 = ~n255 & ~n256;
  assign n258 = ~n199 & ~n202;
  assign n259 = n257 & ~n258;
  assign n260 = ~n257 & n258;
  assign n261 = ~n259 & ~n260;
  assign n262 = n210 & n261;
  assign n263 = ~n210 & ~n261;
  assign n264 = pi23 & ~n263;
  assign n265 = ~n262 & ~n264;
  assign n266 = ~n255 & ~n259;
  assign n267 = ~pi06 & n161;
  assign n268 = ~n218 & ~n267;
  assign n269 = n160 & n213;
  assign n270 = pi03 & pi14;
  assign n271 = n240 & n270;
  assign n272 = pi02 & pi14;
  assign n273 = pi03 & pi13;
  assign n274 = ~n272 & ~n273;
  assign n275 = ~n271 & ~n274;
  assign n276 = n269 & n275;
  assign n277 = ~n269 & ~n275;
  assign n278 = ~n276 & ~n277;
  assign n279 = pi04 & pi12;
  assign n280 = pi05 & pi11;
  assign n281 = ~n279 & ~n280;
  assign n282 = n279 & n280;
  assign n283 = ~n281 & ~n282;
  assign n284 = pi07 & pi09;
  assign n285 = n283 & n284;
  assign n286 = ~n283 & ~n284;
  assign n287 = ~n285 & ~n286;
  assign n288 = n278 & n287;
  assign n289 = ~n278 & ~n287;
  assign n290 = ~n288 & ~n289;
  assign n291 = ~n268 & n290;
  assign n292 = n268 & ~n290;
  assign n293 = ~n291 & ~n292;
  assign n294 = ~n249 & ~n252;
  assign n295 = ~n242 & ~n247;
  assign n296 = ~n233 & ~n236;
  assign n297 = pi06 & pi15;
  assign n298 = n33 & n297;
  assign n299 = pi01 & pi15;
  assign n300 = pi06 & pi10;
  assign n301 = ~n299 & ~n300;
  assign n302 = ~n298 & ~n301;
  assign n303 = ~n296 & n302;
  assign n304 = n296 & ~n302;
  assign n305 = ~n303 & ~n304;
  assign n306 = n295 & ~n305;
  assign n307 = ~n295 & n305;
  assign n308 = ~n306 & ~n307;
  assign n309 = ~n294 & n308;
  assign n310 = n294 & ~n308;
  assign n311 = ~n309 & ~n310;
  assign n312 = n293 & n311;
  assign n313 = ~n293 & ~n311;
  assign n314 = ~n312 & ~n313;
  assign n315 = ~n225 & ~n229;
  assign n316 = n314 & ~n315;
  assign n317 = ~n314 & n315;
  assign n318 = ~n316 & ~n317;
  assign n319 = ~n266 & n318;
  assign n320 = n266 & ~n318;
  assign n321 = ~n319 & ~n320;
  assign n322 = ~n265 & n321;
  assign n323 = ~n316 & ~n319;
  assign n324 = ~n309 & ~n312;
  assign n325 = ~n288 & ~n291;
  assign n326 = ~n271 & ~n276;
  assign n327 = ~n282 & ~n285;
  assign n328 = n298 & ~n327;
  assign n329 = ~n298 & n327;
  assign n330 = ~n328 & ~n329;
  assign n331 = n326 & ~n330;
  assign n332 = ~n326 & n330;
  assign n333 = ~n331 & ~n332;
  assign n334 = ~n325 & n333;
  assign n335 = n325 & ~n333;
  assign n336 = ~n334 & ~n335;
  assign n337 = ~n303 & ~n307;
  assign n338 = pi02 & pi15;
  assign n339 = ~n270 & ~n338;
  assign n340 = pi03 & pi15;
  assign n341 = n272 & n340;
  assign n342 = ~n339 & ~n341;
  assign n343 = pi04 & pi13;
  assign n344 = n342 & n343;
  assign n345 = ~n342 & ~n343;
  assign n346 = ~n344 & ~n345;
  assign n347 = pi05 & pi12;
  assign n348 = pi06 & pi11;
  assign n349 = ~n347 & ~n348;
  assign n350 = pi06 & pi12;
  assign n351 = n280 & n350;
  assign n352 = ~n349 & ~n351;
  assign n353 = pi07 & pi10;
  assign n354 = n352 & n353;
  assign n355 = ~n352 & ~n353;
  assign n356 = ~n354 & ~n355;
  assign n357 = n346 & n356;
  assign n358 = ~n346 & ~n356;
  assign n359 = ~n357 & ~n358;
  assign n360 = ~n337 & n359;
  assign n361 = n337 & ~n359;
  assign n362 = ~n360 & ~n361;
  assign n363 = n336 & n362;
  assign n364 = ~n336 & ~n362;
  assign n365 = ~n363 & ~n364;
  assign n366 = ~n324 & n365;
  assign n367 = n324 & ~n365;
  assign n368 = ~n366 & ~n367;
  assign n369 = ~n323 & n368;
  assign n370 = n323 & ~n368;
  assign n371 = ~n369 & ~n370;
  assign n372 = n322 & n371;
  assign n373 = ~n366 & ~n369;
  assign n374 = ~n334 & ~n363;
  assign n375 = ~n357 & ~n360;
  assign n376 = ~n341 & ~n344;
  assign n377 = n241 & n348;
  assign n378 = pi07 & pi11;
  assign n379 = ~n350 & ~n378;
  assign n380 = ~n377 & ~n379;
  assign n381 = ~n376 & n380;
  assign n382 = n376 & ~n380;
  assign n383 = ~n381 & ~n382;
  assign n384 = ~n375 & n383;
  assign n385 = n375 & ~n383;
  assign n386 = ~n384 & ~n385;
  assign n387 = ~n328 & ~n332;
  assign n388 = pi04 & pi14;
  assign n389 = n340 & n388;
  assign n390 = ~n340 & ~n388;
  assign n391 = ~n389 & ~n390;
  assign n392 = pi05 & pi13;
  assign n393 = n391 & n392;
  assign n394 = ~n391 & ~n392;
  assign n395 = ~n393 & ~n394;
  assign n396 = ~n351 & ~n354;
  assign n397 = n395 & ~n396;
  assign n398 = ~n395 & n396;
  assign n399 = ~n397 & ~n398;
  assign n400 = ~n387 & n399;
  assign n401 = n387 & ~n399;
  assign n402 = ~n400 & ~n401;
  assign n403 = n386 & n402;
  assign n404 = ~n386 & ~n402;
  assign n405 = ~n403 & ~n404;
  assign n406 = ~n374 & n405;
  assign n407 = n374 & ~n405;
  assign n408 = ~n406 & ~n407;
  assign n409 = ~n373 & n408;
  assign n410 = n373 & ~n408;
  assign n411 = ~n409 & ~n410;
  assign n412 = n372 & n411;
  assign n413 = ~n406 & ~n409;
  assign n414 = ~n384 & ~n403;
  assign n415 = ~n397 & ~n400;
  assign n416 = pi05 & pi15;
  assign n417 = n388 & n416;
  assign n418 = pi04 & pi15;
  assign n419 = pi05 & pi14;
  assign n420 = ~n418 & ~n419;
  assign n421 = ~n417 & ~n420;
  assign n422 = pi06 & pi13;
  assign n423 = n421 & n422;
  assign n424 = ~n421 & ~n422;
  assign n425 = ~n423 & ~n424;
  assign n426 = ~n415 & n425;
  assign n427 = n415 & ~n425;
  assign n428 = ~n426 & ~n427;
  assign n429 = ~n377 & ~n381;
  assign n430 = ~n389 & ~n393;
  assign n431 = n241 & ~n430;
  assign n432 = ~n241 & n430;
  assign n433 = ~n431 & ~n432;
  assign n434 = ~n429 & n433;
  assign n435 = n429 & ~n433;
  assign n436 = ~n434 & ~n435;
  assign n437 = n428 & n436;
  assign n438 = ~n428 & ~n436;
  assign n439 = ~n437 & ~n438;
  assign n440 = ~n414 & n439;
  assign n441 = n414 & ~n439;
  assign n442 = ~n440 & ~n441;
  assign n443 = ~n413 & n442;
  assign n444 = n413 & ~n442;
  assign n445 = ~n443 & ~n444;
  assign n446 = n412 & n445;
  assign n447 = ~n440 & ~n443;
  assign n448 = ~n426 & ~n437;
  assign n449 = ~n431 & ~n434;
  assign n450 = ~n417 & ~n423;
  assign n451 = pi06 & pi14;
  assign n452 = n416 & n451;
  assign n453 = ~n416 & ~n451;
  assign n454 = ~n452 & ~n453;
  assign n455 = pi07 & pi13;
  assign n456 = n454 & n455;
  assign n457 = ~n454 & ~n455;
  assign n458 = ~n456 & ~n457;
  assign n459 = ~n450 & n458;
  assign n460 = n450 & ~n458;
  assign n461 = ~n459 & ~n460;
  assign n462 = ~n449 & n461;
  assign n463 = n449 & ~n461;
  assign n464 = ~n462 & ~n463;
  assign n465 = ~n448 & n464;
  assign n466 = n448 & ~n464;
  assign n467 = ~n465 & ~n466;
  assign n468 = ~n447 & n467;
  assign n469 = n447 & ~n467;
  assign n470 = ~n468 & ~n469;
  assign n471 = n446 & n470;
  assign n472 = ~n465 & ~n468;
  assign n473 = ~n459 & ~n462;
  assign n474 = ~n452 & ~n456;
  assign n475 = pi07 & pi14;
  assign n476 = ~n297 & ~n475;
  assign n477 = n297 & n475;
  assign n478 = ~n476 & ~n477;
  assign n479 = ~n474 & n478;
  assign n480 = n474 & ~n478;
  assign n481 = ~n479 & ~n480;
  assign n482 = ~n473 & n481;
  assign n483 = n473 & ~n481;
  assign n484 = ~n482 & ~n483;
  assign n485 = ~n472 & n484;
  assign n486 = n472 & ~n484;
  assign n487 = ~n485 & ~n486;
  assign n488 = n471 & n487;
  assign n489 = ~n482 & ~n485;
  assign n490 = pi07 & pi15;
  assign n491 = ~n451 & ~n479;
  assign n492 = n490 & ~n491;
  assign n493 = ~n479 & ~n490;
  assign n494 = ~n492 & ~n493;
  assign n495 = ~n489 & n494;
  assign n496 = n489 & ~n494;
  assign n497 = ~n495 & ~n496;
  assign n498 = n488 & n497;
  assign n499 = ~n492 & ~n495;
  assign n500 = ~n498 & n499;
  assign n501 = ~n488 & ~n497;
  assign n502 = ~n498 & ~n501;
  assign n503 = ~n471 & ~n487;
  assign n504 = ~n488 & ~n503;
  assign n505 = ~n446 & ~n470;
  assign n506 = ~n471 & ~n505;
  assign n507 = ~n412 & ~n445;
  assign n508 = ~n446 & ~n507;
  assign n509 = ~n372 & ~n411;
  assign n510 = ~n412 & ~n509;
  assign n511 = ~n322 & ~n371;
  assign n512 = ~n372 & ~n511;
  assign n513 = ~pi23 & ~n262;
  assign n514 = ~n263 & ~n513;
  assign n515 = ~n321 & ~n514;
  assign n516 = ~n322 & ~n515;
  assign n517 = ~n262 & ~n263;
  assign n518 = pi23 & ~n517;
  assign n519 = ~pi23 & n517;
  assign n520 = ~n518 & ~n519;
  assign n521 = ~n205 & ~n208;
  assign n522 = pi22 & ~n521;
  assign n523 = ~pi22 & n521;
  assign n524 = ~n522 & ~n523;
  assign n525 = ~n152 & ~n155;
  assign n526 = pi21 & ~n525;
  assign n527 = ~pi21 & n525;
  assign n528 = ~n526 & ~n527;
  assign n529 = ~n113 & ~n116;
  assign n530 = pi20 & ~n529;
  assign n531 = ~pi20 & n529;
  assign n532 = ~n530 & ~n531;
  assign n533 = ~n76 & ~n79;
  assign n534 = pi19 & ~n533;
  assign n535 = ~pi19 & n533;
  assign n536 = ~n534 & ~n535;
  assign po00 = ~n500;
  assign po01 = n502;
  assign po02 = n504;
  assign po03 = n506;
  assign po04 = n508;
  assign po05 = n510;
  assign po06 = n512;
  assign po07 = n516;
  assign po08 = ~n520;
  assign po09 = ~n524;
  assign po10 = ~n528;
  assign po11 = ~n532;
  assign po12 = ~n536;
  assign po13 = 1'b0;
  assign po14 = 1'b0;
  assign po15 = 1'b0;
endmodule
